library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MON6809 is
    port (
        clock:    in std_logic;
        address:  in std_logic_vector(11 downto 0);
        cs_n:     in std_logic;
        data_out: out std_logic_vector(7 downto 0)
    );
end entity;

architecture rtl of MON6809 is
    -- ROM from $F800 to $FFFF (2048 bytes)
    type rom_type is array(0 to 2047) of std_logic_vector(7 downto 0);
    signal rom : rom_type := (
        X"10", X"CE", X"7F", X"FF", X"CE", X"6F", X"FF", X"86", 
        X"03", X"1F", X"8B", X"BD", X"F8", X"AD", X"BD", X"FA", 
        X"C6", X"8E", X"FE", X"94", X"86", X"01", X"3F", X"86", 
        X"3B", X"BD", X"F8", X"C7", X"8E", X"01", X"00", X"1F", 
        X"10", X"BD", X"FA", X"71", X"BD", X"FA", X"68", X"10", 
        X"8E", X"00", X"08", X"1F", X"10", X"BD", X"FA", X"71", 
        X"BD", X"FA", X"68", X"BD", X"F9", X"E3", X"1F", X"20", 
        X"BD", X"FA", X"71", X"BD", X"FA", X"68", X"1F", X"10", 
        X"BD", X"FA", X"71", X"86", X"3B", X"BD", X"F8", X"C7", 
        X"BD", X"FA", X"C6", X"86", X"02", X"C6", X"80", X"8E", 
        X"02", X"00", X"3F", X"86", X"01", X"8E", X"02", X"00", 
        X"3F", X"BD", X"FB", X"2D", X"BD", X"FB", X"33", X"25", 
        X"EA", X"BD", X"FB", X"82", X"20", X"E5", X"34", X"02", 
        X"84", X"7F", X"B1", X"00", X"0D", X"26", X"0A", X"0C", 
        X"22", X"86", X"01", X"97", X"1E", X"86", X"FF", X"97", 
        X"23", X"0C", X"23", X"35", X"82", X"34", X"02", X"9F", 
        X"20", X"A6", X"84", X"97", X"1F", X"0C", X"1F", X"86", 
        X"01", X"97", X"1E", X"35", X"82", X"0F", X"20", X"0F", 
        X"21", X"0F", X"1F", X"39", X"34", X"16", X"9E", X"20", 
        X"27", X"11", X"D6", X"1E", X"D1", X"1F", X"25", X"0B", 
        X"BD", X"FA", X"68", X"96", X"23", X"A1", X"85", X"26", 
        X"F7", X"0C", X"1E", X"35", X"96", X"34", X"02", X"86", 
        X"7F", X"B7", X"D0", X"12", X"86", X"36", X"B7", X"D0", 
        X"11", X"86", X"26", X"B7", X"D0", X"13", X"BD", X"F8", 
        X"8D", X"0F", X"23", X"0F", X"22", X"35", X"82", X"81", 
        X"09", X"26", X"02", X"20", X"C7", X"8D", X"97", X"34", 
        X"06", X"F6", X"D0", X"12", X"C5", X"80", X"2B", X"F9", 
        X"8A", X"80", X"B7", X"D0", X"12", X"35", X"86", X"B6", 
        X"D0", X"11", X"85", X"80", X"2A", X"F9", X"B6", X"D0", 
        X"10", X"84", X"7F", X"39", X"86", X"2E", X"BD", X"F8", 
        X"C7", X"0F", X"05", X"BD", X"F8", X"DF", X"BD", X"F8", 
        X"C7", X"A7", X"80", X"0C", X"05", X"5A", X"C1", X"01", 
        X"2F", X"04", X"81", X"0D", X"26", X"ED", X"86", X"00", 
        X"A7", X"84", X"39", X"34", X"10", X"BD", X"FB", X"AE", 
        X"EC", X"84", X"BD", X"F9", X"C8", X"25", X"02", X"1C", 
        X"FE", X"35", X"90", X"34", X"10", X"BD", X"FB", X"AE", 
        X"EC", X"81", X"BD", X"F9", X"C8", X"25", X"0F", X"34", 
        X"02", X"EC", X"81", X"BD", X"F9", X"C8", X"25", X"06", 
        X"1F", X"89", X"35", X"02", X"1C", X"FE", X"35", X"90", 
        X"BD", X"FB", X"75", X"25", X"09", X"DD", X"06", X"BD", 
        X"FB", X"75", X"25", X"02", X"DD", X"08", X"39", X"BD", 
        X"FB", X"33", X"25", X"1A", X"81", X"01", X"27", X"09", 
        X"BD", X"F9", X"0B", X"25", X"16", X"A7", X"A0", X"20", 
        X"EE", X"8D", X"11", X"1F", X"89", X"A6", X"80", X"A7", 
        X"A0", X"5A", X"26", X"F9", X"20", X"E1", X"1C", X"FE", 
        X"10", X"9F", X"0C", X"39", X"34", X"10", X"86", X"FF", 
        X"4C", X"6D", X"80", X"26", X"FB", X"35", X"90", X"34", 
        X"32", X"A6", X"80", X"A1", X"A0", X"26", X"03", X"4D", 
        X"26", X"F7", X"35", X"B2", X"34", X"36", X"BD", X"F9", 
        X"6C", X"1F", X"89", X"A6", X"80", X"A7", X"A0", X"5A", 
        X"26", X"F9", X"35", X"B6", X"34", X"02", X"8D", X"08", 
        X"1F", X"89", X"35", X"02", X"44", X"44", X"44", X"44", 
        X"84", X"0F", X"8B", X"90", X"19", X"89", X"40", X"19", 
        X"39", X"81", X"30", X"2D", X"18", X"81", X"39", X"2E", 
        X"05", X"84", X"0F", X"1C", X"FE", X"39", X"81", X"41", 
        X"2D", X"0B", X"81", X"46", X"2E", X"07", X"80", X"41", 
        X"8B", X"0A", X"1C", X"FE", X"39", X"1A", X"01", X"39", 
        X"BD", X"F9", X"A9", X"34", X"02", X"1F", X"98", X"BD", 
        X"F9", X"A9", X"48", X"48", X"48", X"48", X"1F", X"89", 
        X"35", X"02", X"59", X"49", X"59", X"49", X"59", X"49", 
        X"59", X"49", X"39", X"34", X"37", X"C6", X"0A", X"34", 
        X"04", X"5F", X"4F", X"68", X"65", X"69", X"64", X"59", 
        X"49", X"10", X"A3", X"66", X"25", X"04", X"A3", X"66", 
        X"6C", X"65", X"6A", X"E4", X"26", X"ED", X"ED", X"66", 
        X"32", X"61", X"35", X"B7", X"34", X"16", X"86", X"58", 
        X"BD", X"F8", X"C7", X"86", X"3D", X"BD", X"F8", X"C7", 
        X"1F", X"10", X"BD", X"FA", X"71", X"35", X"96", X"34", 
        X"36", X"34", X"01", X"86", X"43", X"BD", X"F8", X"C7", 
        X"86", X"43", X"BD", X"F8", X"C7", X"86", X"3D", X"BD", 
        X"F8", X"C7", X"8E", X"FE", X"09", X"10", X"8E", X"00", 
        X"08", X"35", X"04", X"A6", X"80", X"59", X"25", X"02", 
        X"86", X"2D", X"BD", X"F8", X"C7", X"31", X"3F", X"26", 
        X"F2", X"35", X"B6", X"34", X"06", X"1E", X"89", X"86", 
        X"41", X"BD", X"F8", X"C7", X"86", X"3D", X"BD", X"F8", 
        X"C7", X"1E", X"89", X"BD", X"FA", X"7D", X"35", X"86", 
        X"34", X"06", X"1F", X"98", X"BD", X"FA", X"7D", X"35", 
        X"86", X"34", X"06", X"BD", X"FA", X"71", X"35", X"86", 
        X"34", X"06", X"86", X"20", X"BD", X"F8", X"C7", X"35", 
        X"86", X"34", X"06", X"BD", X"FA", X"7D", X"1F", X"98", 
        X"BD", X"FA", X"7D", X"35", X"86", X"34", X"06", X"17", 
        X"FF", X"12", X"17", X"FE", X"42", X"1F", X"98", X"17", 
        X"FE", X"3D", X"35", X"86", X"34", X"06", X"1F", X"89", 
        X"86", X"2E", X"17", X"FE", X"32", X"1F", X"98", X"17", 
        X"FE", X"2D", X"17", X"FF", X"CB", X"35", X"86", X"34", 
        X"16", X"8E", X"02", X"00", X"1F", X"10", X"BD", X"FA", 
        X"71", X"86", X"3A", X"BD", X"F8", X"C7", X"BD", X"FA", 
        X"68", X"5F", X"A6", X"80", X"5C", X"D1", X"05", X"27", 
        X"08", X"BD", X"FA", X"7D", X"BD", X"FA", X"68", X"20", 
        X"F1", X"BD", X"FA", X"C6", X"35", X"16", X"34", X"06", 
        X"86", X"0D", X"BD", X"F8", X"C7", X"35", X"86", X"34", 
        X"12", X"A6", X"80", X"27", X"05", X"BD", X"F8", X"C7", 
        X"20", X"F7", X"35", X"92", X"34", X"06", X"DC", X"06", 
        X"BD", X"FA", X"71", X"35", X"86", X"34", X"36", X"10", 
        X"8E", X"FB", X"23", X"A6", X"80", X"27", X"22", X"81", 
        X"25", X"26", X"19", X"A6", X"80", X"5F", X"6D", X"A5", 
        X"27", X"1B", X"A1", X"A5", X"27", X"03", X"5C", X"20", 
        X"F5", X"8E", X"FB", X"27", X"58", X"10", X"AE", X"A5", 
        X"AD", X"A4", X"20", X"DF", X"17", X"FD", X"B8", X"20", 
        X"DA", X"1C", X"FE", X"35", X"96", X"1A", X"01", X"35", 
        X"96", X"86", X"25", X"16", X"FD", X"A9", X"DC", X"24", 
        X"16", X"FF", X"AC", X"82", X"25", X"6D", X"CD", X"FB", 
        X"19", X"FB", X"1E", X"FB", X"1E", X"8E", X"02", X"00", 
        X"9F", X"00", X"39", X"34", X"24", X"9E", X"00", X"86", 
        X"00", X"97", X"04", X"A6", X"80", X"27", X"22", X"81", 
        X"22", X"27", X"22", X"81", X"20", X"2F", X"F4", X"1F", 
        X"12", X"31", X"3F", X"A6", X"80", X"81", X"20", X"2E", 
        X"FA", X"6F", X"82", X"30", X"01", X"9F", X"00", X"1F", 
        X"21", X"9F", X"02", X"96", X"04", X"1C", X"FE", X"35", 
        X"A4", X"1A", X"01", X"35", X"A4", X"86", X"01", X"97", 
        X"04", X"1F", X"12", X"A6", X"80", X"27", X"E2", X"81", 
        X"22", X"27", X"DE", X"20", X"F6", X"BD", X"FB", X"33", 
        X"25", X"07", X"BD", X"F9", X"1B", X"25", X"02", X"1C", 
        X"FE", X"39", X"10", X"8E", X"FE", X"24", X"BD", X"FB", 
        X"AE", X"6D", X"A4", X"27", X"14", X"9E", X"02", X"BD", 
        X"F9", X"77", X"27", X"05", X"BD", X"FB", X"A4", X"20", 
        X"F0", X"BD", X"FB", X"A4", X"10", X"AE", X"3E", X"6E", 
        X"A4", X"1A", X"01", X"39", X"1F", X"21", X"BD", X"F9", 
        X"6C", X"31", X"A6", X"31", X"23", X"39", X"34", X"16", 
        X"5F", X"A6", X"80", X"27", X"15", X"81", X"22", X"27", 
        X"11", X"81", X"61", X"25", X"08", X"81", X"7B", X"24", 
        X"04", X"80", X"20", X"A7", X"1F", X"5C", X"D1", X"05", 
        X"23", X"E7", X"35", X"96", X"0F", X"1C", X"0F", X"1D", 
        X"0F", X"1B", X"0A", X"1B", X"39", X"0F", X"1B", X"39", 
        X"0D", X"1B", X"27", X"0B", X"34", X"06", X"1F", X"89", 
        X"4F", X"D3", X"1C", X"DD", X"1C", X"35", X"06", X"39", 
        X"4F", X"3F", X"81", X"01", X"26", X"04", X"17", X"FE", 
        X"DE", X"3B", X"81", X"02", X"26", X"04", X"17", X"FC", 
        X"F3", X"3B", X"34", X"02", X"8E", X"FE", X"7C", X"17", 
        X"FE", X"CD", X"35", X"02", X"17", X"FE", X"76", X"17", 
        X"FE", X"BC", X"3B", X"8E", X"FE", X"6A", X"17", X"FE", 
        X"BE", X"3B", X"8E", X"FE", X"73", X"17", X"FE", X"B7", 
        X"3B", X"8E", X"FE", X"51", X"17", X"FE", X"B0", X"3B", 
        X"8E", X"FE", X"59", X"17", X"FE", X"A9", X"3B", X"8E", 
        X"FE", X"49", X"17", X"FE", X"A2", X"3B", X"BD", X"F9", 
        X"38", X"25", X"23", X"10", X"9E", X"06", X"86", X"3A", 
        X"BD", X"FA", X"8C", X"1F", X"20", X"BD", X"FA", X"71", 
        X"BD", X"FA", X"68", X"34", X"20", X"8D", X"12", X"35", 
        X"20", X"8D", X"1C", X"BD", X"FA", X"C6", X"10", X"9C", 
        X"08", X"23", X"E3", X"1C", X"FE", X"39", X"1A", X"01", 
        X"39", X"C6", X"08", X"A6", X"A0", X"BD", X"FA", X"7D", 
        X"BD", X"FA", X"68", X"5A", X"26", X"F5", X"39", X"C6", 
        X"08", X"A6", X"A0", X"81", X"20", X"2C", X"02", X"86", 
        X"2E", X"BD", X"F8", X"C7", X"5A", X"26", X"F2", X"39", 
        X"BD", X"FB", X"75", X"1F", X"02", X"BD", X"F9", X"47", 
        X"25", X"02", X"1C", X"FE", X"39", X"BD", X"FB", X"33", 
        X"25", X"09", X"BD", X"F9", X"1B", X"25", X"F5", X"1F", 
        X"01", X"AD", X"84", X"39", X"BD", X"F9", X"38", X"25", 
        X"45", X"10", X"8E", X"02", X"80", X"BD", X"F9", X"47", 
        X"25", X"3C", X"9E", X"06", X"30", X"1F", X"9F", X"06", 
        X"C6", X"08", X"9E", X"06", X"30", X"01", X"9F", X"06", 
        X"10", X"8E", X"02", X"80", X"9C", X"08", X"24", X"1D", 
        X"A6", X"80", X"A1", X"A0", X"26", X"EC", X"9C", X"08", 
        X"24", X"13", X"10", X"9C", X"0C", X"25", X"E3", X"BD", 
        X"FA", X"DC", X"BD", X"FA", X"68", X"5A", X"26", X"DA", 
        X"BD", X"FA", X"C6", X"20", X"D3", X"C1", X"08", X"27", 
        X"03", X"BD", X"FA", X"C6", X"1C", X"FE", X"39", X"BD", 
        X"F9", X"38", X"25", X"20", X"10", X"8E", X"02", X"80", 
        X"BD", X"F9", X"47", X"25", X"17", X"9E", X"06", X"10", 
        X"8E", X"02", X"80", X"A6", X"A0", X"A7", X"80", X"9C", 
        X"08", X"22", X"07", X"10", X"9C", X"0C", X"25", X"F3", 
        X"20", X"ED", X"1C", X"FE", X"39", X"0F", X"10", X"BD", 
        X"FB", X"75", X"25", X"32", X"DD", X"06", X"BD", X"FB", 
        X"75", X"25", X"2B", X"93", X"06", X"DD", X"0E", X"BD", 
        X"FB", X"75", X"25", X"22", X"DD", X"08", X"9E", X"06", 
        X"10", X"9E", X"08", X"9C", X"08", X"27", X"15", X"22", 
        X"0E", X"0A", X"10", X"1F", X"10", X"D3", X"0E", X"1F", 
        X"01", X"1F", X"20", X"D3", X"0E", X"1F", X"02", X"DC", 
        X"0E", X"BD", X"FD", X"3F", X"1C", X"FE", X"39", X"34", 
        X"36", X"34", X"02", X"A6", X"84", X"A7", X"A4", X"0D", 
        X"10", X"26", X"06", X"30", X"01", X"31", X"21", X"20", 
        X"04", X"30", X"1F", X"31", X"3F", X"35", X"02", X"83", 
        X"00", X"01", X"2A", X"E5", X"1C", X"FE", X"35", X"B6", 
        X"BD", X"FB", X"75", X"25", X"4E", X"DD", X"06", X"BD", 
        X"FB", X"75", X"25", X"47", X"93", X"06", X"DD", X"0E", 
        X"BD", X"FB", X"75", X"25", X"3E", X"DD", X"08", X"9E", 
        X"06", X"10", X"9E", X"08", X"9C", X"08", X"27", X"31", 
        X"86", X"08", X"97", X"11", X"DC", X"0E", X"34", X"06", 
        X"A6", X"80", X"A1", X"A0", X"27", X"13", X"1F", X"10", 
        X"BD", X"FA", X"71", X"BD", X"FA", X"68", X"0A", X"11", 
        X"2A", X"07", X"BD", X"FA", X"C6", X"86", X"08", X"97", 
        X"11", X"35", X"06", X"83", X"00", X"01", X"2A", X"DE", 
        X"96", X"11", X"81", X"08", X"27", X"03", X"BD", X"FA", 
        X"C6", X"1C", X"FE", X"39", X"0F", X"14", X"BD", X"FB", 
        X"75", X"25", X"04", X"DD", X"18", X"0A", X"14", X"BD", 
        X"F8", X"EC", X"0F", X"1A", X"BD", X"FD", X"ED", X"25", 
        X"03", X"1C", X"FE", X"39", X"39", X"86", X"01", X"20", 
        X"16", X"86", X"02", X"20", X"12", X"86", X"03", X"20", 
        X"0E", X"86", X"04", X"20", X"0A", X"86", X"05", X"20", 
        X"06", X"86", X"06", X"20", X"02", X"86", X"07", X"1A", 
        X"01", X"39", X"39", X"39", X"39", X"34", X"14", X"D6", 
        X"1A", X"8E", X"02", X"00", X"A6", X"85", X"27", X"0B", 
        X"5C", X"D7", X"1A", X"C1", X"80", X"27", X"04", X"1C", 
        X"FE", X"35", X"94", X"1A", X"01", X"35", X"94", X"34", 
        X"00", X"45", X"46", X"48", X"49", X"4E", X"5A", X"56", 
        X"C3", X"BA", X"FD", X"EA", X"D3", X"FD", X"EB", X"BB", 
        X"FD", X"EC", X"00", X"48", X"45", X"58", X"53", X"31", 
        X"39", X"4D", X"4F", X"53", X"43", X"00", X"FD", X"60", 
        X"46", X"00", X"FC", X"DF", X"47", X"00", X"FC", X"85", 
        X"48", X"00", X"FC", X"94", X"4C", X"00", X"FD", X"B4", 
        X"4D", X"00", X"FC", X"2E", X"54", X"00", X"FD", X"05", 
        X"3A", X"00", X"FC", X"78", X"58", X"00", X"FB", X"E8", 
        X"00", X"2A", X"4E", X"4D", X"49", X"2A", X"0D", X"0A", 
        X"00", X"2A", X"49", X"52", X"51", X"2A", X"0D", X"0A", 
        X"00", X"2A", X"46", X"49", X"52", X"51", X"2A", X"0D", 
        X"0A", X"00", X"2A", X"53", X"57", X"49", X"2A", X"0D", 
        X"0A", X"00", X"2A", X"53", X"57", X"49", X"32", X"2A", 
        X"0D", X"0A", X"00", X"2A", X"53", X"57", X"49", X"33", 
        X"2A", X"0D", X"0A", X"00", X"55", X"6E", X"64", X"65", 
        X"66", X"69", X"6E", X"65", X"64", X"20", X"73", X"79", 
        X"73", X"74", X"65", X"6D", X"20", X"63", X"61", X"6C", 
        X"6C", X"20", X"24", X"00", X"52", X"45", X"50", X"4C", 
        X"49", X"43", X"41", X"20", X"31", X"20", X"36", X"38", 
        X"30", X"39", X"20", X"4D", X"4F", X"4E", X"49", X"54", 
        X"4F", X"52", X"0D", X"0A", X"00", X"45", X"58", X"49", 
        X"54", X"49", X"4E", X"47", X"2E", X"2E", X"2E", X"0D", 
        X"0A", X"00", X"44", X"55", X"4D", X"50", X"49", X"4E", 
        X"47", X"2E", X"2E", X"2E", X"0D", X"0A", X"00", X"FE", 
        X"D7", X"FE", X"D9", X"FE", X"EC", X"FE", X"FE", X"FF", 
        X"13", X"FF", X"26", X"FF", X"3B", X"FF", X"51", X"4F", 
        X"4B", X"42", X"41", X"44", X"20", X"48", X"45", X"58", 
        X"20", X"52", X"45", X"43", X"4F", X"52", X"44", X"20", 
        X"54", X"59", X"50", X"45", X"4E", X"4F", X"20", X"48", 
        X"45", X"58", X"20", X"52", X"45", X"43", X"4F", X"52", 
        X"44", X"20", X"54", X"59", X"50", X"45", X"42", X"41", 
        X"44", X"20", X"25", X"4D", X"20", X"52", X"45", X"43", 
        X"4F", X"52", X"44", X"20", X"41", X"44", X"44", X"52", 
        X"45", X"53", X"53", X"4E", X"4F", X"20", X"25", X"4D", 
        X"20", X"52", X"45", X"43", X"4F", X"52", X"44", X"20", 
        X"4C", X"45", X"4E", X"47", X"54", X"48", X"4E", X"4F", 
        X"20", X"25", X"4D", X"20", X"52", X"45", X"43", X"4F", 
        X"52", X"44", X"20", X"43", X"48", X"45", X"43", X"4B", 
        X"53", X"55", X"4D", X"42", X"41", X"44", X"20", X"25", 
        X"4D", X"20", X"52", X"45", X"43", X"4F", X"52", X"44", 
        X"20", X"43", X"48", X"45", X"43", X"4B", X"53", X"55", 
        X"4D", X"42", X"41", X"44", X"20", X"25", X"4D", X"20", 
        X"52", X"45", X"43", X"4F", X"52", X"44", X"20", X"44", 
        X"41", X"54", X"41", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"00", X"00", X"FC", X"12", X"FC", X"0B", X"FC", X"20", 
        X"FC", X"19", X"FB", X"EA", X"00", X"F8", X"F8", X"00"
    );
begin
    process(clock)
    begin
        if rising_edge(clock) then
            if cs_n = '0' then
                data_out <= rom(to_integer(unsigned(address)));
            end if;
        end if;
    end process;
end rtl;
