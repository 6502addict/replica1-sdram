library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity BASIC is
    port (
        clock:    in std_logic;
        cs_n:     in std_logic;
        address:  in std_logic_vector(13 downto 0);
        data_out: out std_logic_vector(7 downto 0)
    );
end entity;

architecture rtl of BASIC is
    -- ROM from $E000 to $FFFF (8192 bytes)
    type rom_type is array(0 to 8191) of std_logic_vector(7 downto 0);
    signal rom : rom_type := (
        X"4C", X"A5", X"FC", X"4C", X"EA", X"E2", X"CD", X"E6", 
        X"DB", X"E5", X"A8", X"EA", X"90", X"E7", X"63", X"E9", 
        X"61", X"ED", X"93", X"E9", X"40", X"FD", X"66", X"E7", 
        X"49", X"FD", X"69", X"FD", X"8E", X"FD", X"DB", X"FD", 
        X"41", X"E8", X"39", X"E7", X"0D", X"E7", X"C4", X"E7", 
        X"A6", X"E6", X"1C", X"E7", X"66", X"E7", X"D7", X"E7", 
        X"CB", X"E6", X"E7", X"E7", X"40", X"F4", X"D0", X"E8", 
        X"F3", X"E6", X"2B", X"E5", X"F0", X"E4", X"52", X"E9", 
        X"CF", X"E4", X"55", X"FE", X"BE", X"FE", X"CA", X"FE", 
        X"3D", X"FE", X"35", X"F8", X"C5", X"F8", X"54", X"F8", 
        X"5C", X"F0", X"2D", X"FB", X"4C", X"FC", X"EB", X"F5", 
        X"A8", X"FB", X"2A", X"F4", X"9C", X"F3", X"8B", X"F0", 
        X"CD", X"F3", X"AB", X"F3", X"0C", X"F3", X"20", X"F3", 
        X"4C", X"F3", X"57", X"F3", X"79", X"6A", X"F4", X"79", 
        X"53", X"F4", X"7B", X"2B", X"F6", X"7B", X"0D", X"F7", 
        X"7D", X"36", X"FB", X"50", X"E6", X"EC", X"46", X"E0", 
        X"EC", X"7F", X"6E", X"FB", X"7F", X"47", X"EC", X"64", 
        X"F6", X"EC", X"45", X"4E", X"C4", X"46", X"4F", X"D2", 
        X"4E", X"45", X"58", X"D4", X"44", X"41", X"54", X"C1", 
        X"49", X"4E", X"50", X"55", X"D4", X"44", X"49", X"CD", 
        X"52", X"45", X"41", X"C4", X"43", X"41", X"4C", X"CC", 
        X"50", X"4F", X"D0", X"48", X"49", X"4D", X"45", X"4D", 
        X"BA", X"4C", X"4F", X"4D", X"45", X"4D", X"BA", X"4F", 
        X"4E", X"45", X"52", X"D2", X"52", X"45", X"53", X"55", 
        X"4D", X"C5", X"4C", X"45", X"D4", X"47", X"4F", X"54", 
        X"CF", X"52", X"55", X"CE", X"49", X"C6", X"52", X"45", 
        X"53", X"54", X"4F", X"52", X"C5", X"47", X"4F", X"53", 
        X"55", X"C2", X"52", X"45", X"54", X"55", X"52", X"CE", 
        X"52", X"45", X"CD", X"53", X"54", X"4F", X"D0", X"4F", 
        X"CE", X"50", X"4F", X"4B", X"C5", X"50", X"52", X"49", 
        X"4E", X"D4", X"43", X"4F", X"4E", X"D4", X"4C", X"49", 
        X"53", X"D4", X"43", X"4C", X"45", X"41", X"D2", X"47", 
        X"45", X"D4", X"4E", X"45", X"D7", X"4D", X"45", X"4E", 
        X"D5", X"53", X"41", X"56", X"C5", X"4C", X"4F", X"41", 
        X"C4", X"43", X"4C", X"D3", X"54", X"CF", X"53", X"50", 
        X"43", X"A8", X"54", X"48", X"45", X"CE", X"4E", X"4F", 
        X"D4", X"53", X"54", X"45", X"D0", X"AB", X"AD", X"AA", 
        X"AF", X"DE", X"41", X"4E", X"C4", X"4F", X"D2", X"BE", 
        X"BD", X"BC", X"53", X"47", X"CE", X"49", X"4E", X"D4", 
        X"41", X"42", X"D3", X"46", X"52", X"C5", X"53", X"51", 
        X"D2", X"52", X"4E", X"C4", X"4C", X"4F", X"C7", X"45", 
        X"58", X"D0", X"50", X"45", X"45", X"CB", X"4C", X"45", 
        X"CE", X"53", X"54", X"52", X"A4", X"56", X"41", X"CC", 
        X"41", X"53", X"C3", X"43", X"48", X"52", X"A4", X"4C", 
        X"45", X"46", X"54", X"A4", X"52", X"49", X"47", X"48", 
        X"54", X"A4", X"4D", X"49", X"44", X"A4", X"00", X"4E", 
        X"4F", X"20", X"46", X"4F", X"D2", X"53", X"59", X"4E", 
        X"54", X"41", X"D8", X"4E", X"4F", X"20", X"47", X"4F", 
        X"53", X"55", X"C2", X"4F", X"55", X"54", X"20", X"4F", 
        X"46", X"20", X"44", X"41", X"54", X"C1", X"49", X"4C", 
        X"4C", X"45", X"47", X"20", X"51", X"54", X"D9", X"4F", 
        X"56", X"45", X"52", X"46", X"4C", X"4F", X"D7", X"4F", 
        X"55", X"54", X"20", X"4F", X"46", X"20", X"4D", X"45", 
        X"CD", X"55", X"4E", X"44", X"45", X"46", X"20", X"4C", 
        X"49", X"4E", X"C5", X"42", X"41", X"44", X"20", X"53", 
        X"55", X"42", X"53", X"43", X"D2", X"52", X"45", X"44", 
        X"49", X"CD", X"44", X"49", X"56", X"20", X"42", X"59", 
        X"20", X"B0", X"4E", X"4F", X"54", X"20", X"44", X"49", 
        X"52", X"45", X"43", X"D4", X"57", X"52", X"4F", X"4E", 
        X"47", X"20", X"54", X"59", X"D0", X"4C", X"4F", X"4E", 
        X"47", X"20", X"53", X"54", X"D2", X"4C", X"4F", X"4E", 
        X"47", X"20", X"46", X"4F", X"52", X"4D", X"55", X"4C", 
        X"C1", X"43", X"41", X"4E", X"27", X"54", X"20", X"43", 
        X"4F", X"4E", X"D4", X"4E", X"4F", X"20", X"43", X"46", 
        X"46", X"C1", X"20", X"45", X"52", X"52", X"00", X"20", 
        X"49", X"4E", X"20", X"00", X"0D", X"42", X"52", X"45", 
        X"41", X"4B", X"00", X"BA", X"E8", X"E8", X"E8", X"E8", 
        X"BD", X"01", X"01", X"C9", X"81", X"D0", X"21", X"A5", 
        X"86", X"D0", X"0A", X"BD", X"02", X"01", X"85", X"85", 
        X"BD", X"03", X"01", X"85", X"86", X"DD", X"03", X"01", 
        X"D0", X"07", X"A5", X"85", X"DD", X"02", X"01", X"F0", 
        X"07", X"8A", X"18", X"69", X"12", X"AA", X"D0", X"D8", 
        X"60", X"20", X"91", X"E2", X"85", X"6D", X"84", X"6E", 
        X"38", X"A5", X"96", X"E5", X"9B", X"85", X"5E", X"A8", 
        X"A5", X"97", X"E5", X"9C", X"AA", X"E8", X"98", X"F0", 
        X"23", X"A5", X"96", X"38", X"E5", X"5E", X"85", X"96", 
        X"B0", X"03", X"C6", X"97", X"38", X"A5", X"94", X"E5", 
        X"5E", X"85", X"94", X"B0", X"08", X"C6", X"95", X"90", 
        X"04", X"B1", X"96", X"91", X"94", X"88", X"D0", X"F9", 
        X"B1", X"96", X"91", X"94", X"C6", X"97", X"C6", X"95", 
        X"CA", X"D0", X"F2", X"60", X"0A", X"69", X"36", X"B0", 
        X"35", X"85", X"5E", X"BA", X"E4", X"5E", X"90", X"2E", 
        X"60", X"C4", X"70", X"90", X"28", X"D0", X"04", X"C5", 
        X"6F", X"90", X"22", X"48", X"A2", X"09", X"98", X"48", 
        X"B5", X"93", X"CA", X"10", X"FA", X"20", X"4A", X"F1", 
        X"A2", X"F7", X"68", X"95", X"9D", X"E8", X"30", X"FA", 
        X"68", X"A8", X"68", X"C4", X"70", X"90", X"06", X"D0", 
        X"05", X"C5", X"6F", X"B0", X"01", X"60", X"A2", X"30", 
        X"24", X"D8", X"10", X"03", X"4C", X"AD", X"FD", X"20", 
        X"34", X"FE", X"20", X"31", X"FE", X"BD", X"6F", X"E1", 
        X"48", X"20", X"36", X"FE", X"E8", X"68", X"10", X"F5", 
        X"20", X"0A", X"E5", X"A9", X"02", X"A0", X"E2", X"20", 
        X"0E", X"E9", X"A4", X"76", X"C8", X"F0", X"03", X"20", 
        X"B9", X"F9", X"20", X"34", X"FE", X"A2", X"DD", X"20", 
        X"DC", X"E3", X"86", X"B8", X"84", X"B9", X"46", X"D8", 
        X"20", X"B1", X"00", X"AA", X"F0", X"EC", X"A2", X"FF", 
        X"86", X"76", X"90", X"06", X"20", X"F1", X"E3", X"4C", 
        X"7B", X"E6", X"A6", X"AF", X"86", X"69", X"A6", X"B0", 
        X"86", X"6A", X"20", X"08", X"E8", X"20", X"F1", X"E3", 
        X"84", X"0F", X"20", X"A1", X"E4", X"90", X"44", X"A0", 
        X"01", X"B1", X"9B", X"85", X"5F", X"A5", X"69", X"85", 
        X"5E", X"A5", X"9C", X"85", X"61", X"A5", X"9B", X"88", 
        X"F1", X"9B", X"18", X"65", X"69", X"85", X"69", X"85", 
        X"60", X"A5", X"6A", X"69", X"FF", X"85", X"6A", X"E5", 
        X"9C", X"AA", X"38", X"A5", X"9B", X"E5", X"69", X"A8", 
        X"B0", X"03", X"E8", X"C6", X"61", X"18", X"65", X"5E", 
        X"90", X"03", X"C6", X"5F", X"18", X"B1", X"5E", X"91", 
        X"60", X"C8", X"D0", X"F9", X"E6", X"5F", X"E6", X"61", 
        X"CA", X"D0", X"F2", X"AD", X"00", X"02", X"F0", X"38", 
        X"A5", X"73", X"A4", X"74", X"85", X"6F", X"84", X"70", 
        X"A5", X"69", X"85", X"96", X"65", X"0F", X"85", X"94", 
        X"A4", X"6A", X"84", X"97", X"90", X"01", X"C8", X"84", 
        X"95", X"20", X"41", X"E2", X"A5", X"50", X"A4", X"51", 
        X"8D", X"FE", X"01", X"8C", X"FF", X"01", X"A5", X"6D", 
        X"A4", X"6E", X"85", X"69", X"84", X"6A", X"A4", X"0F", 
        X"B9", X"FB", X"01", X"88", X"91", X"9B", X"D0", X"F8", 
        X"20", X"EC", X"E4", X"A5", X"67", X"A4", X"68", X"85", 
        X"5E", X"84", X"5F", X"18", X"A0", X"01", X"B1", X"5E", 
        X"D0", X"0B", X"A5", X"69", X"85", X"AF", X"A5", X"6A", 
        X"85", X"B0", X"4C", X"EA", X"E2", X"A0", X"04", X"C8", 
        X"B1", X"5E", X"D0", X"FB", X"C8", X"98", X"65", X"5E", 
        X"AA", X"A0", X"00", X"91", X"5E", X"A5", X"5F", X"69", 
        X"00", X"C8", X"91", X"5E", X"86", X"5E", X"85", X"5F", 
        X"90", X"D2", X"A2", X"80", X"86", X"33", X"20", X"11", 
        X"FE", X"E0", X"EF", X"90", X"02", X"A2", X"EF", X"A9", 
        X"00", X"9D", X"00", X"02", X"A2", X"FF", X"A0", X"01", 
        X"60", X"A6", X"B8", X"CA", X"A0", X"04", X"84", X"13", 
        X"24", X"D6", X"10", X"08", X"68", X"68", X"20", X"EC", 
        X"E4", X"4C", X"48", X"E6", X"E8", X"BD", X"00", X"02", 
        X"24", X"13", X"70", X"04", X"C9", X"20", X"F0", X"F4", 
        X"85", X"0E", X"C9", X"22", X"F0", X"63", X"70", X"3C", 
        X"C9", X"3F", X"D0", X"04", X"A9", X"98", X"D0", X"34", 
        X"C9", X"30", X"90", X"04", X"C9", X"3C", X"90", X"2C", 
        X"84", X"AD", X"A9", X"8A", X"85", X"9D", X"A9", X"DF", 
        X"85", X"9E", X"A0", X"00", X"84", X"0F", X"88", X"86", 
        X"B8", X"CA", X"C8", X"D0", X"02", X"E6", X"9E", X"E8", 
        X"BD", X"00", X"02", X"C9", X"20", X"F0", X"F8", X"38", 
        X"F1", X"9D", X"F0", X"EE", X"C9", X"80", X"D0", X"30", 
        X"05", X"0F", X"A4", X"AD", X"E8", X"C8", X"99", X"FB", 
        X"01", X"B9", X"FB", X"01", X"F0", X"39", X"38", X"E9", 
        X"3A", X"F0", X"04", X"C9", X"49", X"D0", X"02", X"85", 
        X"13", X"38", X"E9", X"5A", X"D0", X"97", X"85", X"0E", 
        X"BD", X"00", X"02", X"F0", X"DF", X"C5", X"0E", X"F0", 
        X"DB", X"C8", X"99", X"FB", X"01", X"E8", X"D0", X"F0", 
        X"A6", X"B8", X"E6", X"0F", X"B1", X"9D", X"C8", X"D0", 
        X"02", X"E6", X"9E", X"0A", X"90", X"F6", X"B1", X"9D", 
        X"D0", X"AE", X"BD", X"00", X"02", X"10", X"BB", X"99", 
        X"FD", X"01", X"C6", X"B9", X"A9", X"FF", X"85", X"B8", 
        X"60", X"A5", X"67", X"A6", X"68", X"A0", X"01", X"85", 
        X"9B", X"86", X"9C", X"B1", X"9B", X"F0", X"1F", X"C8", 
        X"C8", X"A5", X"51", X"D1", X"9B", X"90", X"18", X"F0", 
        X"03", X"88", X"D0", X"09", X"A5", X"50", X"88", X"D1", 
        X"9B", X"90", X"0C", X"F0", X"0A", X"88", X"B1", X"9B", 
        X"AA", X"88", X"B1", X"9B", X"B0", X"D7", X"18", X"60", 
        X"D0", X"FD", X"A9", X"00", X"85", X"D6", X"A8", X"91", 
        X"67", X"C8", X"91", X"67", X"A5", X"67", X"69", X"02", 
        X"85", X"69", X"85", X"AF", X"A5", X"68", X"69", X"00", 
        X"85", X"6A", X"85", X"B0", X"20", X"1E", X"E5", X"A9", 
        X"00", X"D0", X"2A", X"A5", X"73", X"A4", X"74", X"85", 
        X"6F", X"84", X"70", X"A5", X"69", X"A4", X"6A", X"85", 
        X"6B", X"84", X"6C", X"85", X"6D", X"84", X"6E", X"20", 
        X"A7", X"E6", X"A2", X"55", X"86", X"52", X"68", X"A8", 
        X"68", X"A2", X"F8", X"9A", X"48", X"98", X"48", X"A9", 
        X"00", X"85", X"7A", X"85", X"14", X"60", X"18", X"A5", 
        X"67", X"69", X"FF", X"85", X"B8", X"A5", X"68", X"69", 
        X"FF", X"85", X"B9", X"60", X"90", X"0A", X"F0", X"08", 
        X"C9", X"A8", X"F0", X"04", X"C9", X"2C", X"D0", X"E5", 
        X"20", X"08", X"E8", X"20", X"A1", X"E4", X"20", X"B7", 
        X"00", X"F0", X"10", X"C9", X"A8", X"F0", X"04", X"C9", 
        X"2C", X"D0", X"84", X"20", X"B1", X"00", X"20", X"08", 
        X"E8", X"D0", X"CA", X"68", X"68", X"A5", X"50", X"05", 
        X"51", X"D0", X"06", X"A9", X"FF", X"85", X"50", X"85", 
        X"51", X"A0", X"01", X"B1", X"9B", X"F0", X"37", X"20", 
        X"B6", X"E6", X"20", X"34", X"FE", X"C8", X"B1", X"9B", 
        X"AA", X"C8", X"B1", X"9B", X"C5", X"51", X"D0", X"04", 
        X"E4", X"50", X"F0", X"02", X"B0", X"20", X"84", X"85", 
        X"20", X"C4", X"F9", X"A9", X"20", X"A4", X"85", X"29", 
        X"7F", X"20", X"36", X"FE", X"C8", X"B1", X"9B", X"D0", 
        X"1B", X"A8", X"B1", X"9B", X"AA", X"C8", X"B1", X"9B", 
        X"86", X"9B", X"85", X"9C", X"D0", X"C3", X"20", X"34", 
        X"FE", X"4C", X"48", X"E6", X"C8", X"D0", X"02", X"E6", 
        X"9E", X"B1", X"9D", X"60", X"10", X"DB", X"38", X"E9", 
        X"7F", X"AA", X"84", X"85", X"A0", X"8A", X"84", X"9D", 
        X"A0", X"DF", X"84", X"9E", X"A0", X"FF", X"CA", X"F0", 
        X"07", X"20", X"A4", X"E5", X"10", X"FB", X"30", X"F6", 
        X"20", X"2E", X"FE", X"20", X"A4", X"E5", X"30", X"05", 
        X"20", X"36", X"FE", X"D0", X"F6", X"20", X"36", X"FE", 
        X"A9", X"20", X"D0", X"A9", X"A9", X"80", X"85", X"14", 
        X"20", X"42", X"E8", X"20", X"13", X"E2", X"D0", X"05", 
        X"8A", X"69", X"0F", X"AA", X"9A", X"68", X"68", X"A9", 
        X"09", X"20", X"84", X"E2", X"20", X"9F", X"E7", X"18", 
        X"98", X"65", X"B8", X"48", X"A5", X"B9", X"69", X"00", 
        X"48", X"A5", X"76", X"48", X"A5", X"75", X"48", X"A9", 
        X"A2", X"20", X"69", X"EC", X"20", X"1A", X"EB", X"20", 
        X"17", X"EB", X"A5", X"A2", X"09", X"7F", X"25", X"9E", 
        X"85", X"9E", X"A9", X"25", X"A0", X"E6", X"85", X"5E", 
        X"84", X"5F", X"4C", X"D0", X"EB", X"A9", X"BD", X"A0", 
        X"F5", X"20", X"9E", X"F7", X"20", X"B7", X"00", X"C9", 
        X"A6", X"D0", X"06", X"20", X"B1", X"00", X"20", X"17", 
        X"EB", X"20", X"27", X"F8", X"20", X"C5", X"EB", X"A5", 
        X"86", X"48", X"A5", X"85", X"48", X"A9", X"81", X"48", 
        X"BA", X"86", X"F8", X"20", X"B6", X"E6", X"A5", X"B8", 
        X"A4", X"B9", X"A6", X"76", X"E8", X"F0", X"04", X"85", 
        X"79", X"84", X"7A", X"A0", X"00", X"B1", X"B8", X"D0", 
        X"3F", X"A0", X"02", X"B1", X"B8", X"18", X"F0", X"1C", 
        X"C8", X"B1", X"B8", X"85", X"75", X"C8", X"B1", X"B8", 
        X"85", X"76", X"98", X"65", X"B8", X"85", X"B8", X"90", 
        X"02", X"E6", X"B9", X"20", X"B1", X"00", X"20", X"86", 
        X"E6", X"4C", X"48", X"E6", X"F0", X"62", X"F0", X"2D", 
        X"E9", X"80", X"90", X"11", X"C9", X"40", X"B0", X"14", 
        X"0A", X"A8", X"B9", X"07", X"E0", X"48", X"B9", X"06", 
        X"E0", X"48", X"4C", X"B1", X"00", X"4C", X"42", X"E8", 
        X"C9", X"3A", X"F0", X"D7", X"4C", X"72", X"EC", X"38", 
        X"A5", X"67", X"E9", X"01", X"A4", X"68", X"B0", X"01", 
        X"88", X"85", X"7D", X"84", X"7E", X"60", X"AD", X"10", 
        X"D0", X"C9", X"83", X"F0", X"01", X"60", X"20", X"F2", 
        X"FD", X"A2", X"FF", X"24", X"D8", X"10", X"03", X"4C", 
        X"AD", X"FD", X"C9", X"03", X"B0", X"01", X"18", X"D0", 
        X"3C", X"A5", X"B8", X"A4", X"B9", X"A6", X"76", X"E8", 
        X"F0", X"0C", X"85", X"79", X"84", X"7A", X"A5", X"75", 
        X"A4", X"76", X"85", X"77", X"84", X"78", X"68", X"68", 
        X"A9", X"0C", X"A0", X"E2", X"90", X"03", X"4C", X"DF", 
        X"E2", X"4C", X"EA", X"E2", X"D0", X"17", X"A2", X"82", 
        X"A4", X"7A", X"D0", X"03", X"4C", X"C0", X"E2", X"A5", 
        X"79", X"85", X"B8", X"84", X"B9", X"A5", X"77", X"A4", 
        X"78", X"85", X"75", X"84", X"76", X"60", X"08", X"C6", 
        X"76", X"28", X"D0", X"03", X"4C", X"EC", X"E4", X"20", 
        X"F3", X"E4", X"4C", X"31", X"E7", X"A9", X"03", X"20", 
        X"84", X"E2", X"A5", X"B9", X"48", X"A5", X"B8", X"48", 
        X"A5", X"76", X"48", X"A5", X"75", X"48", X"A9", X"92", 
        X"48", X"20", X"B7", X"00", X"20", X"3A", X"E7", X"4C", 
        X"48", X"E6", X"20", X"08", X"E8", X"20", X"A2", X"E7", 
        X"A5", X"76", X"C5", X"51", X"B0", X"0B", X"98", X"38", 
        X"65", X"B8", X"A6", X"B9", X"90", X"07", X"E8", X"B0", 
        X"04", X"A5", X"67", X"A6", X"68", X"20", X"A5", X"E4", 
        X"90", X"1E", X"A5", X"9B", X"E9", X"01", X"85", X"B8", 
        X"A5", X"9C", X"E9", X"00", X"85", X"B9", X"60", X"D0", 
        X"FD", X"A9", X"FF", X"85", X"85", X"20", X"13", X"E2", 
        X"9A", X"C9", X"92", X"F0", X"0B", X"A2", X"0C", X"2C", 
        X"A2", X"3A", X"4C", X"C0", X"E2", X"4C", X"72", X"EC", 
        X"68", X"68", X"C0", X"10", X"F0", X"3B", X"85", X"75", 
        X"68", X"85", X"76", X"68", X"85", X"B8", X"68", X"85", 
        X"B9", X"20", X"9F", X"E7", X"98", X"18", X"65", X"B8", 
        X"85", X"B8", X"90", X"02", X"E6", X"B9", X"60", X"A2", 
        X"3A", X"2C", X"A2", X"00", X"86", X"0D", X"A0", X"00", 
        X"84", X"0E", X"A5", X"0E", X"A6", X"0D", X"85", X"0D", 
        X"86", X"0E", X"B1", X"B8", X"F0", X"E8", X"C5", X"0E", 
        X"F0", X"E4", X"C8", X"C9", X"22", X"D0", X"F3", X"F0", 
        X"E9", X"68", X"68", X"68", X"60", X"20", X"2B", X"EB", 
        X"20", X"B7", X"00", X"C9", X"8E", X"F0", X"05", X"A9", 
        X"A4", X"20", X"69", X"EC", X"A5", X"9D", X"D0", X"05", 
        X"20", X"A2", X"E7", X"F0", X"B7", X"20", X"B7", X"00", 
        X"B0", X"03", X"4C", X"3A", X"E7", X"4C", X"86", X"E6", 
        X"20", X"BE", X"F3", X"48", X"C9", X"92", X"F0", X"04", 
        X"C9", X"8E", X"D0", X"89", X"C6", X"A1", X"D0", X"04", 
        X"68", X"4C", X"88", X"E6", X"20", X"B1", X"00", X"20", 
        X"08", X"E8", X"C9", X"2C", X"F0", X"EE", X"68", X"60", 
        X"A2", X"00", X"86", X"50", X"86", X"51", X"B0", X"F7", 
        X"E9", X"2F", X"85", X"0D", X"A5", X"51", X"85", X"5E", 
        X"C9", X"19", X"B0", X"D4", X"A5", X"50", X"0A", X"26", 
        X"5E", X"0A", X"26", X"5E", X"65", X"50", X"85", X"50", 
        X"A5", X"5E", X"65", X"51", X"85", X"51", X"06", X"50", 
        X"26", X"51", X"A5", X"50", X"65", X"0D", X"85", X"50", 
        X"90", X"02", X"E6", X"51", X"20", X"B1", X"00", X"4C", 
        X"0E", X"E8", X"20", X"6C", X"ED", X"85", X"85", X"84", 
        X"86", X"A9", X"AF", X"20", X"69", X"EC", X"A5", X"12", 
        X"48", X"A5", X"11", X"48", X"20", X"2B", X"EB", X"68", 
        X"2A", X"20", X"1D", X"EB", X"D0", X"18", X"68", X"10", 
        X"12", X"20", X"17", X"F8", X"20", X"8B", X"EE", X"A0", 
        X"00", X"A5", X"A0", X"91", X"85", X"C8", X"A5", X"A1", 
        X"91", X"85", X"60", X"4C", X"CC", X"F7", X"68", X"A0", 
        X"02", X"B1", X"A0", X"C5", X"70", X"90", X"17", X"D0", 
        X"07", X"88", X"B1", X"A0", X"C5", X"6F", X"90", X"0E", 
        X"A4", X"A1", X"C4", X"6A", X"90", X"08", X"D0", X"0D", 
        X"A5", X"A0", X"C5", X"69", X"B0", X"07", X"A5", X"A0", 
        X"A4", X"A1", X"4C", X"B3", X"E8", X"A0", X"00", X"B1", 
        X"A0", X"20", X"9B", X"F0", X"A5", X"8C", X"A4", X"8D", 
        X"85", X"AB", X"84", X"AC", X"20", X"9A", X"F2", X"A9", 
        X"9D", X"A0", X"00", X"85", X"8C", X"84", X"8D", X"20", 
        X"FB", X"F2", X"A0", X"00", X"B1", X"8C", X"91", X"85", 
        X"C8", X"B1", X"8C", X"91", X"85", X"C8", X"B1", X"8C", 
        X"91", X"85", X"60", X"20", X"11", X"E9", X"20", X"B7", 
        X"00", X"F0", X"1F", X"F0", X"F5", X"C9", X"A3", X"18", 
        X"F0", X"1B", X"C9", X"2C", X"F0", X"25", X"C9", X"3B", 
        X"F0", X"21", X"20", X"2B", X"EB", X"24", X"11", X"30", 
        X"E2", X"20", X"D4", X"F9", X"20", X"AD", X"F0", X"4C", 
        X"CB", X"E8", X"4C", X"34", X"FE", X"20", X"BB", X"F3", 
        X"C9", X"29", X"F0", X"03", X"4C", X"72", X"EC", X"E8", 
        X"CA", X"D0", X"06", X"20", X"B1", X"00", X"4C", X"D3", 
        X"E8", X"20", X"2E", X"FE", X"D0", X"F2", X"20", X"AD", 
        X"F0", X"20", X"C6", X"F2", X"AA", X"A0", X"00", X"E8", 
        X"CA", X"F0", X"AF", X"B1", X"5E", X"20", X"36", X"FE", 
        X"C8", X"4C", X"18", X"E9", X"A5", X"15", X"F0", X"12", 
        X"30", X"04", X"A0", X"FF", X"D0", X"04", X"A5", X"7B", 
        X"A4", X"7C", X"85", X"75", X"84", X"76", X"4C", X"72", 
        X"EC", X"68", X"24", X"D8", X"10", X"05", X"A2", X"FE", 
        X"4C", X"AD", X"FD", X"A9", X"9F", X"A0", X"EA", X"20", 
        X"0E", X"E9", X"A5", X"79", X"A4", X"7A", X"85", X"B8", 
        X"84", X"B9", X"60", X"20", X"81", X"F0", X"A2", X"01", 
        X"A0", X"02", X"A9", X"00", X"8D", X"01", X"02", X"A9", 
        X"40", X"4C", X"9D", X"E9", X"C9", X"22", X"D0", X"0E", 
        X"20", X"31", X"EC", X"A9", X"3B", X"20", X"69", X"EC", 
        X"20", X"11", X"E9", X"4C", X"79", X"E9", X"20", X"31", 
        X"FE", X"20", X"81", X"F0", X"A9", X"2C", X"8D", X"FF", 
        X"01", X"20", X"DA", X"E3", X"AD", X"00", X"02", X"C9", 
        X"03", X"D0", X"10", X"4C", X"C1", X"E6", X"20", X"31", 
        X"FE", X"4C", X"DA", X"E3", X"A6", X"7D", X"A4", X"7E", 
        X"A9", X"98", X"2C", X"A9", X"00", X"85", X"15", X"86", 
        X"7F", X"84", X"80", X"20", X"6C", X"ED", X"85", X"85", 
        X"84", X"86", X"A5", X"B8", X"A4", X"B9", X"85", X"87", 
        X"84", X"88", X"A6", X"7F", X"A4", X"80", X"86", X"B8", 
        X"84", X"B9", X"20", X"B7", X"00", X"D0", X"1C", X"24", 
        X"15", X"50", X"0C", X"20", X"F2", X"FD", X"8D", X"00", 
        X"02", X"A2", X"FF", X"A0", X"01", X"D0", X"08", X"30", 
        X"7F", X"20", X"31", X"FE", X"20", X"8E", X"E9", X"86", 
        X"B8", X"84", X"B9", X"20", X"B1", X"00", X"24", X"11", 
        X"10", X"31", X"24", X"15", X"50", X"09", X"E8", X"86", 
        X"B8", X"A9", X"00", X"85", X"0D", X"F0", X"0C", X"85", 
        X"0D", X"C9", X"22", X"F0", X"07", X"A9", X"3A", X"85", 
        X"0D", X"A9", X"2C", X"18", X"85", X"0E", X"A5", X"B8", 
        X"A4", X"B9", X"69", X"00", X"90", X"01", X"C8", X"20", 
        X"B3", X"F0", X"20", X"03", X"F4", X"20", X"77", X"E8", 
        X"4C", X"22", X"EA", X"48", X"AD", X"00", X"02", X"F0", 
        X"30", X"68", X"20", X"EC", X"F8", X"A5", X"12", X"20", 
        X"5F", X"E8", X"20", X"B7", X"00", X"F0", X"07", X"C9", 
        X"2C", X"F0", X"03", X"4C", X"24", X"E9", X"A5", X"B8", 
        X"A4", X"B9", X"85", X"7F", X"84", X"80", X"A5", X"87", 
        X"A4", X"88", X"85", X"B8", X"84", X"B9", X"20", X"B7", 
        X"00", X"F0", X"33", X"20", X"67", X"EC", X"4C", X"A3", 
        X"E9", X"A5", X"15", X"D0", X"CC", X"4C", X"39", X"E9", 
        X"20", X"9F", X"E7", X"C8", X"AA", X"D0", X"12", X"A2", 
        X"14", X"C8", X"B1", X"B8", X"F0", X"5F", X"C8", X"B1", 
        X"B8", X"85", X"7B", X"C8", X"B1", X"B8", X"C8", X"85", 
        X"7C", X"B1", X"B8", X"AA", X"20", X"94", X"E7", X"E0", 
        X"83", X"D0", X"DD", X"4C", X"DB", X"E9", X"A5", X"7F", 
        X"A4", X"80", X"A6", X"15", X"10", X"03", X"4C", X"B1", 
        X"E6", X"A0", X"00", X"B1", X"7F", X"F0", X"07", X"A9", 
        X"8F", X"A0", X"EA", X"4C", X"0E", X"E9", X"60", X"3F", 
        X"45", X"58", X"54", X"52", X"41", X"20", X"49", X"47", 
        X"4E", X"4F", X"52", X"45", X"44", X"0D", X"00", X"3F", 
        X"52", X"45", X"45", X"4E", X"54", X"45", X"52", X"0D", 
        X"00", X"D0", X"04", X"A0", X"00", X"F0", X"03", X"20", 
        X"6C", X"ED", X"85", X"85", X"84", X"86", X"20", X"13", 
        X"E2", X"F0", X"04", X"A2", X"00", X"F0", X"69", X"9A", 
        X"E8", X"E8", X"E8", X"E8", X"8A", X"E8", X"E8", X"E8", 
        X"E8", X"E8", X"E8", X"86", X"60", X"A0", X"01", X"20", 
        X"9E", X"F7", X"BA", X"BD", X"09", X"01", X"85", X"A2", 
        X"A5", X"85", X"A4", X"86", X"20", X"68", X"F4", X"20", 
        X"CC", X"F7", X"A0", X"01", X"20", X"59", X"F8", X"BA", 
        X"38", X"FD", X"09", X"01", X"F0", X"17", X"BD", X"0F", 
        X"01", X"85", X"75", X"BD", X"10", X"01", X"85", X"76", 
        X"BD", X"12", X"01", X"85", X"B8", X"BD", X"11", X"01", 
        X"85", X"B9", X"4C", X"48", X"E6", X"8A", X"69", X"11", 
        X"AA", X"9A", X"20", X"B7", X"00", X"C9", X"2C", X"D0", 
        X"F1", X"20", X"B1", X"00", X"20", X"AF", X"EA", X"20", 
        X"2B", X"EB", X"18", X"24", X"38", X"24", X"11", X"30", 
        X"03", X"B0", X"03", X"60", X"B0", X"FD", X"A2", X"65", 
        X"4C", X"C0", X"E2", X"A6", X"B8", X"D0", X"02", X"C6", 
        X"B9", X"C6", X"B8", X"A2", X"00", X"24", X"48", X"8A", 
        X"48", X"A9", X"01", X"20", X"84", X"E2", X"20", X"10", 
        X"EC", X"A9", X"00", X"85", X"89", X"20", X"B7", X"00", 
        X"38", X"E9", X"AE", X"90", X"17", X"C9", X"03", X"B0", 
        X"13", X"C9", X"01", X"2A", X"49", X"01", X"45", X"89", 
        X"C5", X"89", X"90", X"61", X"85", X"89", X"20", X"B1", 
        X"00", X"4C", X"48", X"EB", X"A6", X"89", X"D0", X"2C", 
        X"B0", X"7B", X"69", X"07", X"90", X"77", X"65", X"11", 
        X"D0", X"03", X"4C", X"5D", X"F2", X"69", X"FF", X"85", 
        X"5E", X"0A", X"65", X"5E", X"A8", X"68", X"D9", X"6C", 
        X"E0", X"B0", X"67", X"20", X"1A", X"EB", X"48", X"20", 
        X"AD", X"EB", X"68", X"A4", X"87", X"10", X"17", X"AA", 
        X"F0", X"56", X"D0", X"5F", X"46", X"11", X"8A", X"2A", 
        X"A6", X"B8", X"D0", X"02", X"C6", X"B9", X"C6", X"B8", 
        X"A0", X"1B", X"85", X"89", X"D0", X"D7", X"D9", X"6C", 
        X"E0", X"B0", X"48", X"90", X"D9", X"B9", X"6E", X"E0", 
        X"48", X"B9", X"6D", X"E0", X"48", X"20", X"C0", X"EB", 
        X"A5", X"89", X"4C", X"36", X"EB", X"4C", X"72", X"EC", 
        X"A5", X"A2", X"BE", X"6C", X"E0", X"A8", X"68", X"85", 
        X"5E", X"E6", X"5E", X"68", X"85", X"5F", X"98", X"48", 
        X"20", X"17", X"F8", X"A5", X"A1", X"48", X"A5", X"A0", 
        X"48", X"A5", X"9F", X"48", X"A5", X"9E", X"48", X"A5", 
        X"9D", X"48", X"6C", X"5E", X"00", X"A0", X"FF", X"68", 
        X"F0", X"23", X"C9", X"64", X"F0", X"03", X"20", X"1A", 
        X"EB", X"84", X"87", X"68", X"4A", X"85", X"16", X"68", 
        X"85", X"A5", X"68", X"85", X"A6", X"68", X"85", X"A7", 
        X"68", X"85", X"A8", X"68", X"85", X"A9", X"68", X"85", 
        X"AA", X"45", X"A2", X"85", X"AB", X"A5", X"9D", X"60", 
        X"A9", X"00", X"85", X"11", X"20", X"B1", X"00", X"B0", 
        X"03", X"4C", X"EC", X"F8", X"20", X"FC", X"ED", X"B0", 
        X"5D", X"C9", X"2E", X"F0", X"F4", X"C9", X"A8", X"F0", 
        X"4E", X"C9", X"A7", X"F0", X"E7", X"C9", X"22", X"D0", 
        X"0F", X"A5", X"B8", X"A4", X"B9", X"69", X"00", X"90", 
        X"01", X"C8", X"20", X"AD", X"F0", X"4C", X"03", X"F4", 
        X"C9", X"A5", X"D0", X"10", X"A0", X"18", X"D0", X"31", 
        X"A5", X"9D", X"D0", X"03", X"A0", X"01", X"2C", X"A0", 
        X"00", X"4C", X"7D", X"F0", X"C9", X"B1", X"90", X"03", 
        X"4C", X"A2", X"EC", X"20", X"64", X"EC", X"20", X"2B", 
        X"EB", X"A9", X"29", X"2C", X"A9", X"28", X"2C", X"A9", 
        X"2C", X"A0", X"00", X"D1", X"B8", X"D0", X"03", X"4C", 
        X"B1", X"00", X"A2", X"06", X"4C", X"C0", X"E2", X"A0", 
        X"15", X"68", X"68", X"4C", X"87", X"EB", X"20", X"6C", 
        X"ED", X"85", X"A0", X"84", X"A1", X"A6", X"11", X"F0", 
        X"05", X"A2", X"00", X"86", X"AC", X"60", X"A6", X"12", 
        X"10", X"0D", X"A0", X"00", X"B1", X"A0", X"AA", X"C8", 
        X"B1", X"A0", X"A8", X"8A", X"4C", X"70", X"F0", X"4C", 
        X"9E", X"F7", X"0A", X"48", X"AA", X"20", X"B1", X"00", 
        X"E0", X"7D", X"90", X"20", X"20", X"64", X"EC", X"20", 
        X"2B", X"EB", X"20", X"67", X"EC", X"20", X"1C", X"EB", 
        X"68", X"AA", X"A5", X"A1", X"48", X"A5", X"A0", X"48", 
        X"8A", X"48", X"20", X"BE", X"F3", X"68", X"A8", X"8A", 
        X"48", X"4C", X"D1", X"EC", X"20", X"5B", X"EC", X"68", 
        X"A8", X"B9", X"E8", X"DF", X"85", X"91", X"B9", X"E9", 
        X"DF", X"85", X"92", X"20", X"90", X"00", X"4C", X"1A", 
        X"EB", X"A5", X"A5", X"05", X"9D", X"D0", X"0B", X"A5", 
        X"A5", X"F0", X"04", X"A5", X"9D", X"D0", X"03", X"A0", 
        X"00", X"2C", X"A0", X"01", X"4C", X"7D", X"F0", X"20", 
        X"1D", X"EB", X"B0", X"13", X"A5", X"AA", X"09", X"7F", 
        X"25", X"A6", X"85", X"A6", X"A9", X"A5", X"A0", X"00", 
        X"20", X"57", X"F8", X"AA", X"4C", X"42", X"ED", X"A9", 
        X"00", X"85", X"11", X"C6", X"89", X"20", X"C6", X"F2", 
        X"85", X"9D", X"86", X"9E", X"84", X"9F", X"A5", X"A8", 
        X"A4", X"A9", X"20", X"CA", X"F2", X"86", X"A8", X"84", 
        X"A9", X"AA", X"38", X"E5", X"9D", X"F0", X"08", X"A9", 
        X"01", X"90", X"04", X"A6", X"9D", X"A9", X"FF", X"85", 
        X"A2", X"A0", X"FF", X"E8", X"C8", X"CA", X"D0", X"07", 
        X"A6", X"A2", X"30", X"0F", X"18", X"90", X"0C", X"B1", 
        X"A8", X"D1", X"9E", X"F0", X"EF", X"A2", X"FF", X"B0", 
        X"02", X"A2", X"01", X"E8", X"8A", X"2A", X"25", X"16", 
        X"F0", X"02", X"A9", X"01", X"4C", X"38", X"F8", X"20", 
        X"67", X"EC", X"AA", X"20", X"71", X"ED", X"20", X"B7", 
        X"00", X"D0", X"F4", X"60", X"A2", X"00", X"20", X"B7", 
        X"00", X"86", X"10", X"85", X"81", X"20", X"B7", X"00", 
        X"20", X"FC", X"ED", X"B0", X"03", X"4C", X"72", X"EC", 
        X"A2", X"00", X"86", X"11", X"86", X"12", X"20", X"B1", 
        X"00", X"90", X"05", X"20", X"FC", X"ED", X"90", X"0B", 
        X"AA", X"20", X"B1", X"00", X"90", X"FB", X"20", X"FC", 
        X"ED", X"B0", X"F6", X"C9", X"24", X"D0", X"06", X"A9", 
        X"FF", X"85", X"11", X"D0", X"10", X"C9", X"25", X"D0", 
        X"13", X"A5", X"14", X"30", X"D0", X"A9", X"80", X"85", 
        X"12", X"05", X"81", X"85", X"81", X"8A", X"09", X"80", 
        X"AA", X"20", X"B1", X"00", X"86", X"82", X"38", X"05", 
        X"14", X"E9", X"28", X"D0", X"03", X"4C", X"9D", X"EE", 
        X"24", X"14", X"30", X"02", X"70", X"F7", X"A9", X"00", 
        X"85", X"14", X"A5", X"69", X"A6", X"6A", X"A0", X"00", 
        X"86", X"9C", X"85", X"9B", X"E4", X"6C", X"D0", X"04", 
        X"C5", X"6B", X"F0", X"21", X"A5", X"81", X"D1", X"9B", 
        X"D0", X"08", X"A5", X"82", X"C8", X"D1", X"9B", X"F0", 
        X"6B", X"88", X"18", X"A5", X"9B", X"69", X"07", X"90", 
        X"E1", X"E8", X"D0", X"DC", X"C9", X"5B", X"B0", X"03", 
        X"C9", X"41", X"60", X"18", X"60", X"68", X"48", X"C9", 
        X"80", X"D0", X"0F", X"BA", X"BD", X"02", X"01", X"C9", 
        X"EC", X"D0", X"07", X"A9", X"18", X"A0", X"EE", X"60", 
        X"00", X"00", X"A5", X"6B", X"A4", X"6C", X"85", X"9B", 
        X"84", X"9C", X"A5", X"6D", X"A4", X"6E", X"85", X"96", 
        X"84", X"97", X"18", X"69", X"07", X"90", X"01", X"C8", 
        X"85", X"94", X"84", X"95", X"20", X"41", X"E2", X"A5", 
        X"94", X"A4", X"95", X"C8", X"85", X"6B", X"84", X"6C", 
        X"A0", X"00", X"A5", X"81", X"91", X"9B", X"C8", X"A5", 
        X"82", X"91", X"9B", X"A9", X"00", X"C8", X"91", X"9B", 
        X"C8", X"91", X"9B", X"C8", X"91", X"9B", X"C8", X"91", 
        X"9B", X"C8", X"91", X"9B", X"A5", X"9B", X"18", X"69", 
        X"02", X"A4", X"9C", X"90", X"01", X"C8", X"85", X"83", 
        X"84", X"84", X"60", X"A5", X"0F", X"0A", X"69", X"05", 
        X"65", X"9B", X"A4", X"9C", X"90", X"01", X"C8", X"85", 
        X"94", X"84", X"95", X"60", X"90", X"80", X"00", X"00", 
        X"00", X"20", X"B1", X"00", X"20", X"17", X"EB", X"A5", 
        X"A2", X"30", X"0D", X"A5", X"9D", X"C9", X"90", X"90", 
        X"09", X"A9", X"7C", X"A0", X"EE", X"20", X"57", X"F8", 
        X"D0", X"7E", X"4C", X"94", X"F8", X"A5", X"14", X"D0", 
        X"47", X"A5", X"10", X"05", X"12", X"48", X"A5", X"11", 
        X"48", X"A0", X"00", X"98", X"48", X"A5", X"82", X"48", 
        X"A5", X"81", X"48", X"20", X"81", X"EE", X"68", X"85", 
        X"81", X"68", X"85", X"82", X"68", X"A8", X"BA", X"BD", 
        X"02", X"01", X"48", X"BD", X"01", X"01", X"48", X"A5", 
        X"A0", X"9D", X"02", X"01", X"A5", X"A1", X"9D", X"01", 
        X"01", X"C8", X"20", X"B7", X"00", X"C9", X"2C", X"F0", 
        X"D2", X"84", X"0F", X"20", X"61", X"EC", X"68", X"85", 
        X"11", X"68", X"85", X"12", X"29", X"7F", X"85", X"10", 
        X"A6", X"6B", X"A5", X"6C", X"86", X"9B", X"85", X"9C", 
        X"C5", X"6E", X"D0", X"04", X"E4", X"6D", X"F0", X"3F", 
        X"A0", X"00", X"B1", X"9B", X"C8", X"C5", X"81", X"D0", 
        X"06", X"A5", X"82", X"D1", X"9B", X"F0", X"16", X"C8", 
        X"B1", X"9B", X"18", X"65", X"9B", X"AA", X"C8", X"B1", 
        X"9B", X"65", X"9C", X"90", X"D7", X"A2", X"44", X"2C", 
        X"A2", X"1F", X"4C", X"C0", X"E2", X"A2", X"4E", X"A5", 
        X"10", X"D0", X"F7", X"A5", X"14", X"F0", X"02", X"38", 
        X"60", X"20", X"6B", X"EE", X"A5", X"0F", X"A0", X"04", 
        X"D1", X"9B", X"D0", X"E1", X"4C", X"C9", X"EF", X"A5", 
        X"14", X"F0", X"05", X"A2", X"14", X"4C", X"C0", X"E2", 
        X"20", X"6B", X"EE", X"20", X"91", X"E2", X"A0", X"00", 
        X"84", X"AE", X"A2", X"05", X"A5", X"81", X"91", X"9B", 
        X"10", X"01", X"CA", X"C8", X"A5", X"82", X"91", X"9B", 
        X"10", X"02", X"CA", X"CA", X"86", X"AD", X"A5", X"0F", 
        X"C8", X"C8", X"C8", X"91", X"9B", X"A2", X"0B", X"A9", 
        X"00", X"24", X"10", X"50", X"08", X"68", X"18", X"69", 
        X"01", X"AA", X"68", X"69", X"00", X"C8", X"91", X"9B", 
        X"C8", X"8A", X"91", X"9B", X"20", X"2B", X"F0", X"86", 
        X"AD", X"85", X"AE", X"A4", X"5E", X"C6", X"0F", X"D0", 
        X"DC", X"65", X"95", X"B0", X"5D", X"85", X"95", X"A8", 
        X"8A", X"65", X"94", X"90", X"03", X"C8", X"F0", X"52", 
        X"20", X"91", X"E2", X"85", X"6D", X"84", X"6E", X"A9", 
        X"00", X"E6", X"AE", X"A4", X"AD", X"F0", X"05", X"88", 
        X"91", X"94", X"D0", X"FB", X"C6", X"95", X"C6", X"AE", 
        X"D0", X"F5", X"E6", X"95", X"38", X"A5", X"6D", X"E5", 
        X"9B", X"A0", X"02", X"91", X"9B", X"A5", X"6E", X"C8", 
        X"E5", X"9C", X"91", X"9B", X"A5", X"10", X"D0", X"62", 
        X"C8", X"B1", X"9B", X"85", X"0F", X"A9", X"00", X"85", 
        X"AD", X"85", X"AE", X"C8", X"68", X"AA", X"85", X"A0", 
        X"68", X"85", X"A1", X"D1", X"9B", X"90", X"0E", X"D0", 
        X"06", X"C8", X"8A", X"D1", X"9B", X"90", X"07", X"4C", 
        X"15", X"EF", X"4C", X"BE", X"E2", X"C8", X"A5", X"AE", 
        X"05", X"AD", X"18", X"F0", X"0A", X"20", X"2B", X"F0", 
        X"8A", X"65", X"A0", X"AA", X"98", X"A4", X"5E", X"65", 
        X"A1", X"86", X"AD", X"C6", X"0F", X"D0", X"CA", X"85", 
        X"AE", X"A2", X"05", X"A5", X"81", X"10", X"01", X"CA", 
        X"A5", X"82", X"10", X"02", X"CA", X"CA", X"86", X"64", 
        X"A9", X"00", X"20", X"34", X"F0", X"8A", X"65", X"94", 
        X"85", X"83", X"98", X"65", X"95", X"85", X"84", X"A8", 
        X"A5", X"83", X"60", X"84", X"5E", X"B1", X"9B", X"85", 
        X"64", X"88", X"B1", X"9B", X"85", X"65", X"A9", X"10", 
        X"85", X"99", X"A2", X"00", X"A0", X"00", X"8A", X"0A", 
        X"AA", X"98", X"2A", X"A8", X"B0", X"A4", X"06", X"AD", 
        X"26", X"AE", X"90", X"0B", X"18", X"8A", X"65", X"64", 
        X"AA", X"98", X"65", X"65", X"A8", X"B0", X"93", X"C6", 
        X"99", X"D0", X"E3", X"60", X"A5", X"11", X"F0", X"03", 
        X"20", X"C6", X"F2", X"20", X"4A", X"F1", X"38", X"A5", 
        X"6F", X"E5", X"6D", X"A8", X"A5", X"70", X"E5", X"6E", 
        X"A2", X"00", X"86", X"11", X"85", X"9E", X"84", X"9F", 
        X"A2", X"90", X"4C", X"40", X"F8", X"A9", X"00", X"F0", 
        X"EF", X"A6", X"76", X"E8", X"D0", X"A4", X"A2", X"5B", 
        X"4C", X"C0", X"E2", X"20", X"1A", X"EB", X"A0", X"00", 
        X"20", X"D6", X"F9", X"68", X"68", X"A9", X"FF", X"A0", 
        X"00", X"F0", X"12", X"A6", X"A0", X"A4", X"A1", X"86", 
        X"8C", X"84", X"8D", X"20", X"18", X"F1", X"86", X"9E", 
        X"84", X"9F", X"85", X"9D", X"60", X"A2", X"22", X"86", 
        X"0D", X"86", X"0E", X"85", X"AB", X"84", X"AC", X"85", 
        X"9E", X"84", X"9F", X"A0", X"FF", X"C8", X"B1", X"AB", 
        X"F0", X"0C", X"C5", X"0D", X"F0", X"04", X"C5", X"0E", 
        X"D0", X"F3", X"C9", X"22", X"F0", X"01", X"18", X"84", 
        X"9D", X"98", X"65", X"AB", X"85", X"AD", X"A6", X"AC", 
        X"90", X"01", X"E8", X"86", X"AE", X"A5", X"AC", X"F0", 
        X"04", X"C9", X"02", X"D0", X"0B", X"98", X"20", X"9B", 
        X"F0", X"A6", X"AB", X"A4", X"AC", X"20", X"A8", X"F2", 
        X"A6", X"52", X"E0", X"5E", X"D0", X"05", X"A2", X"76", 
        X"4C", X"C0", X"E2", X"A5", X"9D", X"95", X"00", X"A5", 
        X"9E", X"95", X"01", X"A5", X"9F", X"95", X"02", X"A0", 
        X"00", X"86", X"A0", X"84", X"A1", X"88", X"84", X"11", 
        X"86", X"53", X"E8", X"E8", X"E8", X"86", X"52", X"60", 
        X"46", X"13", X"48", X"49", X"FF", X"38", X"65", X"6F", 
        X"A4", X"70", X"B0", X"01", X"88", X"C4", X"6E", X"90", 
        X"11", X"D0", X"04", X"C5", X"6D", X"90", X"0B", X"85", 
        X"6F", X"84", X"70", X"85", X"71", X"84", X"72", X"AA", 
        X"68", X"60", X"A2", X"30", X"A5", X"13", X"30", X"B8", 
        X"20", X"4A", X"F1", X"A9", X"80", X"85", X"13", X"68", 
        X"D0", X"D0", X"A6", X"73", X"A5", X"74", X"86", X"6F", 
        X"85", X"70", X"A0", X"00", X"84", X"8B", X"A5", X"6D", 
        X"A6", X"6E", X"85", X"9B", X"86", X"9C", X"A9", X"55", 
        X"A2", X"00", X"85", X"5E", X"86", X"5F", X"C5", X"52", 
        X"F0", X"05", X"20", X"E9", X"F1", X"F0", X"F7", X"A9", 
        X"07", X"85", X"8F", X"A5", X"69", X"A6", X"6A", X"85", 
        X"5E", X"86", X"5F", X"E4", X"6C", X"D0", X"04", X"C5", 
        X"6B", X"F0", X"05", X"20", X"DF", X"F1", X"F0", X"F3", 
        X"85", X"94", X"86", X"95", X"A9", X"03", X"85", X"8F", 
        X"A5", X"94", X"A6", X"95", X"E4", X"6E", X"D0", X"07", 
        X"C5", X"6D", X"D0", X"03", X"4C", X"28", X"F2", X"85", 
        X"5E", X"86", X"5F", X"A0", X"00", X"B1", X"5E", X"AA", 
        X"C8", X"B1", X"5E", X"08", X"C8", X"B1", X"5E", X"65", 
        X"94", X"85", X"94", X"C8", X"B1", X"5E", X"65", X"95", 
        X"85", X"95", X"28", X"10", X"D3", X"8A", X"30", X"D0", 
        X"C8", X"B1", X"5E", X"A0", X"00", X"0A", X"69", X"05", 
        X"65", X"5E", X"85", X"5E", X"90", X"02", X"E6", X"5F", 
        X"A6", X"5F", X"E4", X"95", X"D0", X"04", X"C5", X"94", 
        X"F0", X"BA", X"20", X"E9", X"F1", X"F0", X"F3", X"B1", 
        X"5E", X"30", X"35", X"C8", X"B1", X"5E", X"10", X"30", 
        X"C8", X"B1", X"5E", X"F0", X"2B", X"C8", X"B1", X"5E", 
        X"AA", X"C8", X"B1", X"5E", X"C5", X"70", X"90", X"06", 
        X"D0", X"1E", X"E4", X"6F", X"B0", X"1A", X"C5", X"9C", 
        X"90", X"16", X"D0", X"04", X"E4", X"9B", X"90", X"10", 
        X"86", X"9B", X"85", X"9C", X"A5", X"5E", X"A6", X"5F", 
        X"85", X"8A", X"86", X"8B", X"A5", X"8F", X"85", X"91", 
        X"A5", X"8F", X"18", X"65", X"5E", X"85", X"5E", X"90", 
        X"02", X"E6", X"5F", X"A6", X"5F", X"A0", X"00", X"60", 
        X"A6", X"8B", X"F0", X"F7", X"A5", X"91", X"29", X"04", 
        X"4A", X"A8", X"85", X"91", X"B1", X"8A", X"65", X"9B", 
        X"85", X"96", X"A5", X"9C", X"69", X"00", X"85", X"97", 
        X"A5", X"6F", X"A6", X"70", X"85", X"94", X"86", X"95", 
        X"20", X"48", X"E2", X"A4", X"91", X"C8", X"A5", X"94", 
        X"91", X"8A", X"AA", X"E6", X"95", X"A5", X"95", X"C8", 
        X"91", X"8A", X"4C", X"4E", X"F1", X"A5", X"A1", X"48", 
        X"A5", X"A0", X"48", X"20", X"10", X"EC", X"20", X"1C", 
        X"EB", X"68", X"85", X"AB", X"68", X"85", X"AC", X"A0", 
        X"00", X"B1", X"AB", X"18", X"71", X"A0", X"90", X"05", 
        X"A2", X"6E", X"4C", X"C0", X"E2", X"20", X"9B", X"F0", 
        X"20", X"9A", X"F2", X"A5", X"8C", X"A4", X"8D", X"20", 
        X"CA", X"F2", X"20", X"AC", X"F2", X"A5", X"AB", X"A4", 
        X"AC", X"20", X"CA", X"F2", X"20", X"F0", X"F0", X"4C", 
        X"45", X"EB", X"A0", X"00", X"B1", X"AB", X"48", X"C8", 
        X"B1", X"AB", X"AA", X"C8", X"B1", X"AB", X"A8", X"68", 
        X"86", X"5E", X"84", X"5F", X"A8", X"F0", X"0A", X"48", 
        X"88", X"B1", X"5E", X"91", X"71", X"98", X"D0", X"F8", 
        X"68", X"18", X"65", X"71", X"85", X"71", X"90", X"02", 
        X"E6", X"72", X"60", X"20", X"1C", X"EB", X"A5", X"A0", 
        X"A4", X"A1", X"85", X"5E", X"84", X"5F", X"20", X"FB", 
        X"F2", X"08", X"A0", X"00", X"B1", X"5E", X"48", X"C8", 
        X"B1", X"5E", X"AA", X"C8", X"B1", X"5E", X"A8", X"68", 
        X"28", X"D0", X"13", X"C4", X"70", X"D0", X"0F", X"E4", 
        X"6F", X"D0", X"0B", X"48", X"18", X"65", X"6F", X"85", 
        X"6F", X"90", X"02", X"E6", X"70", X"68", X"86", X"5E", 
        X"84", X"5F", X"60", X"C4", X"54", X"D0", X"0C", X"C5", 
        X"53", X"D0", X"08", X"85", X"52", X"E9", X"03", X"85", 
        X"53", X"A0", X"00", X"60", X"20", X"C1", X"F3", X"8A", 
        X"48", X"A9", X"01", X"20", X"A3", X"F0", X"68", X"A0", 
        X"00", X"91", X"9E", X"68", X"68", X"4C", X"F0", X"F0", 
        X"20", X"7F", X"F3", X"D1", X"8C", X"98", X"90", X"04", 
        X"B1", X"8C", X"AA", X"98", X"48", X"8A", X"48", X"20", 
        X"A3", X"F0", X"A5", X"8C", X"A4", X"8D", X"20", X"CA", 
        X"F2", X"68", X"A8", X"68", X"18", X"65", X"5E", X"85", 
        X"5E", X"90", X"02", X"E6", X"5F", X"98", X"20", X"AC", 
        X"F2", X"4C", X"F0", X"F0", X"20", X"7F", X"F3", X"18", 
        X"F1", X"8C", X"49", X"FF", X"4C", X"26", X"F3", X"A9", 
        X"FF", X"85", X"A1", X"20", X"B7", X"00", X"C9", X"29", 
        X"F0", X"06", X"20", X"67", X"EC", X"20", X"BE", X"F3", 
        X"20", X"7F", X"F3", X"CA", X"8A", X"48", X"18", X"A2", 
        X"00", X"F1", X"8C", X"B0", X"B8", X"49", X"FF", X"C5", 
        X"A1", X"90", X"B3", X"A5", X"A1", X"B0", X"AF", X"20", 
        X"61", X"EC", X"68", X"A8", X"68", X"85", X"91", X"68", 
        X"68", X"68", X"AA", X"68", X"85", X"8C", X"68", X"85", 
        X"8D", X"A5", X"91", X"48", X"98", X"48", X"A0", X"00", 
        X"8A", X"F0", X"1D", X"60", X"20", X"A2", X"F3", X"4C", 
        X"7D", X"F0", X"20", X"C3", X"F2", X"A2", X"00", X"86", 
        X"11", X"A8", X"60", X"20", X"A2", X"F3", X"F0", X"08", 
        X"A0", X"00", X"B1", X"5E", X"A8", X"4C", X"7D", X"F0", 
        X"4C", X"18", X"EF", X"20", X"B1", X"00", X"20", X"17", 
        X"EB", X"20", X"87", X"EE", X"A6", X"A0", X"D0", X"F0", 
        X"A6", X"A1", X"4C", X"B7", X"00", X"20", X"A2", X"F3", 
        X"D0", X"03", X"4C", X"F8", X"F4", X"A6", X"B8", X"A4", 
        X"B9", X"86", X"AD", X"84", X"AE", X"A6", X"5E", X"86", 
        X"B8", X"18", X"65", X"5E", X"85", X"60", X"A6", X"5F", 
        X"86", X"B9", X"90", X"01", X"E8", X"86", X"61", X"A0", 
        X"00", X"B1", X"60", X"48", X"A9", X"00", X"91", X"60", 
        X"20", X"B7", X"00", X"20", X"EC", X"F8", X"68", X"A0", 
        X"00", X"91", X"60", X"A6", X"AD", X"A4", X"AE", X"86", 
        X"B8", X"84", X"B9", X"60", X"20", X"17", X"EB", X"20", 
        X"18", X"F4", X"20", X"67", X"EC", X"4C", X"BE", X"F3", 
        X"A5", X"9D", X"C9", X"91", X"B0", X"9A", X"20", X"94", 
        X"F8", X"A5", X"A0", X"A4", X"A1", X"84", X"50", X"85", 
        X"51", X"60", X"A5", X"50", X"48", X"A5", X"51", X"48", 
        X"20", X"18", X"F4", X"A0", X"00", X"B1", X"50", X"A8", 
        X"68", X"85", X"51", X"68", X"85", X"50", X"4C", X"7D", 
        X"F0", X"20", X"0C", X"F4", X"8A", X"A0", X"00", X"91", 
        X"50", X"60", X"A9", X"04", X"A0", X"FB", X"4C", X"68", 
        X"F4", X"20", X"8B", X"F6", X"A5", X"A2", X"49", X"FF", 
        X"85", X"A2", X"45", X"AA", X"85", X"AB", X"A5", X"9D", 
        X"4C", X"6B", X"F4", X"20", X"9A", X"F5", X"90", X"3C", 
        X"20", X"8B", X"F6", X"D0", X"03", X"4C", X"F8", X"F7", 
        X"A6", X"AC", X"86", X"92", X"A2", X"A5", X"A5", X"A5", 
        X"A8", X"F0", X"CE", X"38", X"E5", X"9D", X"F0", X"24", 
        X"90", X"12", X"84", X"9D", X"A4", X"AA", X"84", X"A2", 
        X"49", X"FF", X"69", X"00", X"A0", X"00", X"84", X"92", 
        X"A2", X"9D", X"D0", X"04", X"A0", X"00", X"84", X"AC", 
        X"C9", X"F9", X"30", X"C7", X"A8", X"A5", X"AC", X"56", 
        X"01", X"20", X"B1", X"F5", X"24", X"AB", X"10", X"57", 
        X"A0", X"9D", X"E0", X"A5", X"F0", X"02", X"A0", X"A5", 
        X"38", X"49", X"FF", X"65", X"92", X"85", X"AC", X"B9", 
        X"04", X"00", X"F5", X"04", X"85", X"A1", X"B9", X"03", 
        X"00", X"F5", X"03", X"85", X"A0", X"B9", X"02", X"00", 
        X"F5", X"02", X"85", X"9F", X"B9", X"01", X"00", X"F5", 
        X"01", X"85", X"9E", X"B0", X"03", X"20", X"48", X"F5", 
        X"A0", X"00", X"98", X"18", X"A6", X"9E", X"D0", X"4A", 
        X"A6", X"9F", X"86", X"9E", X"A6", X"A0", X"86", X"9F", 
        X"A6", X"A1", X"86", X"A0", X"A6", X"AC", X"86", X"A1", 
        X"84", X"AC", X"69", X"08", X"C9", X"20", X"D0", X"E4", 
        X"A9", X"00", X"85", X"9D", X"85", X"A2", X"60", X"65", 
        X"92", X"85", X"AC", X"A5", X"A1", X"65", X"A9", X"85", 
        X"A1", X"A5", X"A0", X"65", X"A8", X"85", X"A0", X"A5", 
        X"9F", X"65", X"A7", X"85", X"9F", X"A5", X"9E", X"65", 
        X"A6", X"85", X"9E", X"4C", X"37", X"F5", X"69", X"01", 
        X"06", X"AC", X"26", X"A1", X"26", X"A0", X"26", X"9F", 
        X"26", X"9E", X"10", X"F2", X"38", X"E5", X"9D", X"B0", 
        X"C7", X"49", X"FF", X"69", X"01", X"85", X"9D", X"90", 
        X"0E", X"E6", X"9D", X"F0", X"42", X"66", X"9E", X"66", 
        X"9F", X"66", X"A0", X"66", X"A1", X"66", X"AC", X"60", 
        X"A5", X"A2", X"49", X"FF", X"85", X"A2", X"A5", X"9E", 
        X"49", X"FF", X"85", X"9E", X"A5", X"9F", X"49", X"FF", 
        X"85", X"9F", X"A5", X"A0", X"49", X"FF", X"85", X"A0", 
        X"A5", X"A1", X"49", X"FF", X"85", X"A1", X"A5", X"AC", 
        X"49", X"FF", X"85", X"AC", X"E6", X"AC", X"D0", X"0E", 
        X"E6", X"A1", X"D0", X"0A", X"E6", X"A0", X"D0", X"06", 
        X"E6", X"9F", X"D0", X"02", X"E6", X"9E", X"60", X"A2", 
        X"28", X"4C", X"C0", X"E2", X"A2", X"61", X"B4", X"04", 
        X"84", X"AC", X"B4", X"03", X"94", X"04", X"B4", X"02", 
        X"94", X"03", X"B4", X"01", X"94", X"02", X"A4", X"A4", 
        X"94", X"01", X"69", X"08", X"30", X"E8", X"F0", X"E6", 
        X"E9", X"08", X"A8", X"A5", X"AC", X"B0", X"14", X"16", 
        X"01", X"90", X"02", X"F6", X"01", X"76", X"01", X"76", 
        X"01", X"76", X"02", X"76", X"03", X"76", X"04", X"6A", 
        X"C8", X"D0", X"EC", X"18", X"60", X"81", X"00", X"00", 
        X"00", X"00", X"03", X"7F", X"5E", X"56", X"CB", X"79", 
        X"80", X"13", X"9B", X"0B", X"64", X"80", X"76", X"38", 
        X"93", X"16", X"82", X"38", X"AA", X"3B", X"20", X"80", 
        X"35", X"04", X"F3", X"34", X"81", X"35", X"04", X"F3", 
        X"34", X"80", X"80", X"00", X"00", X"00", X"80", X"31", 
        X"72", X"17", X"F8", X"20", X"27", X"F8", X"F0", X"02", 
        X"10", X"03", X"4C", X"18", X"EF", X"A5", X"9D", X"E9", 
        X"7F", X"48", X"A9", X"80", X"85", X"9D", X"A9", X"D7", 
        X"A0", X"F5", X"20", X"68", X"F4", X"A9", X"DC", X"A0", 
        X"F5", X"20", X"0B", X"F7", X"A9", X"BD", X"A0", X"F5", 
        X"20", X"51", X"F4", X"A9", X"C2", X"A0", X"F5", X"20", 
        X"FA", X"FB", X"A9", X"E1", X"A0", X"F5", X"20", X"68", 
        X"F4", X"68", X"20", X"76", X"F9", X"A9", X"E6", X"A0", 
        X"F5", X"20", X"8B", X"F6", X"D0", X"01", X"60", X"20", 
        X"B6", X"F6", X"A9", X"00", X"85", X"62", X"85", X"63", 
        X"85", X"64", X"85", X"65", X"A5", X"AC", X"20", X"58", 
        X"F6", X"A5", X"A1", X"20", X"58", X"F6", X"A5", X"A0", 
        X"20", X"58", X"F6", X"A5", X"9F", X"20", X"58", X"F6", 
        X"A5", X"9E", X"20", X"5D", X"F6", X"4C", X"8B", X"F7", 
        X"D0", X"03", X"4C", X"84", X"F5", X"4A", X"09", X"80", 
        X"A8", X"90", X"19", X"18", X"A5", X"65", X"65", X"A9", 
        X"85", X"65", X"A5", X"64", X"65", X"A8", X"85", X"64", 
        X"A5", X"63", X"65", X"A7", X"85", X"63", X"A5", X"62", 
        X"65", X"A6", X"85", X"62", X"66", X"62", X"66", X"63", 
        X"66", X"64", X"66", X"65", X"66", X"AC", X"98", X"4A", 
        X"D0", X"D6", X"60", X"85", X"5E", X"84", X"5F", X"A0", 
        X"04", X"B1", X"5E", X"85", X"A9", X"88", X"B1", X"5E", 
        X"85", X"A8", X"88", X"B1", X"5E", X"85", X"A7", X"88", 
        X"B1", X"5E", X"85", X"AA", X"45", X"A2", X"85", X"AB", 
        X"A5", X"AA", X"09", X"80", X"85", X"A6", X"88", X"B1", 
        X"5E", X"85", X"A5", X"A5", X"9D", X"60", X"A5", X"A5", 
        X"F0", X"1C", X"18", X"65", X"9D", X"90", X"04", X"30", 
        X"1A", X"18", X"2C", X"10", X"11", X"69", X"80", X"85", 
        X"9D", X"F0", X"02", X"A5", X"AB", X"85", X"A2", X"60", 
        X"A5", X"A2", X"49", X"FF", X"30", X"05", X"68", X"68", 
        X"4C", X"F8", X"F4", X"4C", X"7F", X"F5", X"20", X"08", 
        X"F8", X"AA", X"F0", X"10", X"18", X"69", X"02", X"B0", 
        X"F2", X"A2", X"00", X"86", X"AB", X"20", X"78", X"F4", 
        X"E6", X"9D", X"F0", X"E7", X"60", X"84", X"20", X"00", 
        X"00", X"00", X"20", X"08", X"F8", X"A9", X"F5", X"A0", 
        X"F6", X"A2", X"00", X"86", X"AB", X"20", X"9E", X"F7", 
        X"4C", X"0E", X"F7", X"20", X"8B", X"F6", X"F0", X"76", 
        X"20", X"17", X"F8", X"A9", X"00", X"38", X"E5", X"9D", 
        X"85", X"9D", X"20", X"B6", X"F6", X"E6", X"9D", X"F0", 
        X"BA", X"A2", X"FC", X"A9", X"01", X"A4", X"A6", X"C4", 
        X"9E", X"D0", X"10", X"A4", X"A7", X"C4", X"9F", X"D0", 
        X"0A", X"A4", X"A8", X"C4", X"A0", X"D0", X"04", X"A4", 
        X"A9", X"C4", X"A1", X"08", X"2A", X"90", X"09", X"E8", 
        X"95", X"65", X"F0", X"32", X"10", X"34", X"A9", X"01", 
        X"28", X"B0", X"0E", X"06", X"A9", X"26", X"A8", X"26", 
        X"A7", X"26", X"A6", X"B0", X"E6", X"30", X"CE", X"10", 
        X"E2", X"A8", X"A5", X"A9", X"E5", X"A1", X"85", X"A9", 
        X"A5", X"A8", X"E5", X"A0", X"85", X"A8", X"A5", X"A7", 
        X"E5", X"9F", X"85", X"A7", X"A5", X"A6", X"E5", X"9E", 
        X"85", X"A6", X"98", X"4C", X"4B", X"F7", X"A9", X"40", 
        X"D0", X"CE", X"0A", X"0A", X"0A", X"0A", X"0A", X"0A", 
        X"85", X"AC", X"28", X"4C", X"8B", X"F7", X"A2", X"53", 
        X"4C", X"C0", X"E2", X"A5", X"62", X"85", X"9E", X"A5", 
        X"63", X"85", X"9F", X"A5", X"64", X"85", X"A0", X"A5", 
        X"65", X"85", X"A1", X"4C", X"D8", X"F4", X"85", X"5E", 
        X"84", X"5F", X"A0", X"04", X"B1", X"5E", X"85", X"A1", 
        X"88", X"B1", X"5E", X"85", X"A0", X"88", X"B1", X"5E", 
        X"85", X"9F", X"88", X"B1", X"5E", X"85", X"A2", X"09", 
        X"80", X"85", X"9E", X"88", X"B1", X"5E", X"85", X"9D", 
        X"84", X"AC", X"60", X"A2", X"98", X"2C", X"A2", X"93", 
        X"A0", X"00", X"F0", X"04", X"A6", X"85", X"A4", X"86", 
        X"20", X"17", X"F8", X"86", X"5E", X"84", X"5F", X"A0", 
        X"04", X"A5", X"A1", X"91", X"5E", X"88", X"A5", X"A0", 
        X"91", X"5E", X"88", X"A5", X"9F", X"91", X"5E", X"88", 
        X"A5", X"A2", X"09", X"7F", X"25", X"9E", X"91", X"5E", 
        X"88", X"A5", X"9D", X"91", X"5E", X"84", X"AC", X"60", 
        X"A5", X"AA", X"85", X"A2", X"A2", X"05", X"B5", X"A4", 
        X"95", X"9C", X"CA", X"D0", X"F9", X"86", X"AC", X"60", 
        X"20", X"17", X"F8", X"A2", X"06", X"B5", X"9C", X"95", 
        X"A4", X"CA", X"D0", X"F9", X"86", X"AC", X"60", X"A5", 
        X"9D", X"F0", X"FB", X"06", X"AC", X"90", X"F7", X"20", 
        X"70", X"F5", X"D0", X"F2", X"4C", X"39", X"F5", X"A5", 
        X"9D", X"F0", X"09", X"A5", X"A2", X"2A", X"A9", X"FF", 
        X"B0", X"02", X"A9", X"01", X"60", X"20", X"27", X"F8", 
        X"85", X"9E", X"A9", X"00", X"85", X"9F", X"A2", X"88", 
        X"A5", X"9E", X"49", X"FF", X"2A", X"A9", X"00", X"85", 
        X"A1", X"85", X"A0", X"86", X"9D", X"85", X"AC", X"85", 
        X"A2", X"4C", X"D3", X"F4", X"46", X"A2", X"60", X"85", 
        X"60", X"84", X"61", X"A0", X"00", X"B1", X"60", X"C8", 
        X"AA", X"F0", X"C4", X"B1", X"60", X"45", X"A2", X"30", 
        X"C2", X"E4", X"9D", X"D0", X"21", X"B1", X"60", X"09", 
        X"80", X"C5", X"9E", X"D0", X"19", X"C8", X"B1", X"60", 
        X"C5", X"9F", X"D0", X"12", X"C8", X"B1", X"60", X"C5", 
        X"A0", X"D0", X"0B", X"C8", X"A9", X"7F", X"C5", X"AC", 
        X"B1", X"60", X"E5", X"A1", X"F0", X"25", X"6A", X"45", 
        X"A2", X"4C", X"2D", X"F8", X"A5", X"9D", X"F0", X"4A", 
        X"38", X"E9", X"A0", X"24", X"A2", X"10", X"09", X"AA", 
        X"A9", X"FF", X"85", X"A4", X"20", X"4E", X"F5", X"8A", 
        X"A2", X"9D", X"C9", X"F9", X"10", X"06", X"20", X"9A", 
        X"F5", X"84", X"A4", X"60", X"A8", X"A5", X"A2", X"29", 
        X"80", X"46", X"9E", X"05", X"9E", X"85", X"9E", X"20", 
        X"B1", X"F5", X"84", X"A4", X"60", X"A5", X"9D", X"C9", 
        X"A0", X"B0", X"20", X"20", X"94", X"F8", X"84", X"AC", 
        X"A5", X"A2", X"84", X"A2", X"49", X"80", X"2A", X"A9", 
        X"A0", X"85", X"9D", X"A5", X"A1", X"85", X"0D", X"4C", 
        X"D3", X"F4", X"85", X"9E", X"85", X"9F", X"85", X"A0", 
        X"85", X"A1", X"A8", X"60", X"A0", X"00", X"A2", X"0A", 
        X"94", X"99", X"CA", X"10", X"FB", X"90", X"0F", X"C9", 
        X"2D", X"D0", X"04", X"86", X"A3", X"F0", X"04", X"C9", 
        X"2B", X"D0", X"05", X"20", X"B1", X"00", X"90", X"5B", 
        X"C9", X"2E", X"F0", X"2E", X"C9", X"45", X"D0", X"30", 
        X"20", X"B1", X"00", X"90", X"17", X"C9", X"A8", X"F0", 
        X"0E", X"C9", X"2D", X"F0", X"0A", X"C9", X"A7", X"F0", 
        X"08", X"C9", X"2B", X"F0", X"04", X"D0", X"07", X"66", 
        X"9C", X"20", X"B1", X"00", X"90", X"5B", X"24", X"9C", 
        X"10", X"0E", X"A9", X"00", X"38", X"E5", X"9A", X"4C", 
        X"42", X"F9", X"66", X"9B", X"24", X"9B", X"50", X"C3", 
        X"A5", X"9A", X"38", X"E5", X"99", X"85", X"9A", X"F0", 
        X"12", X"10", X"09", X"20", X"FA", X"F6", X"E6", X"9A", 
        X"D0", X"F9", X"F0", X"07", X"20", X"DE", X"F6", X"C6", 
        X"9A", X"D0", X"F9", X"A5", X"A3", X"30", X"01", X"60", 
        X"4C", X"6F", X"FB", X"48", X"24", X"9B", X"10", X"02", 
        X"E6", X"99", X"20", X"DE", X"F6", X"68", X"29", X"0F", 
        X"20", X"76", X"F9", X"4C", X"03", X"F9", X"48", X"20", 
        X"08", X"F8", X"68", X"20", X"38", X"F8", X"A5", X"AA", 
        X"45", X"A2", X"85", X"AB", X"A6", X"9D", X"4C", X"6B", 
        X"F4", X"A5", X"9A", X"C9", X"0A", X"90", X"09", X"A9", 
        X"64", X"24", X"9C", X"30", X"10", X"4C", X"7F", X"F5", 
        X"0A", X"0A", X"18", X"65", X"9A", X"0A", X"A0", X"00", 
        X"71", X"B8", X"38", X"E9", X"30", X"85", X"9A", X"4C", 
        X"29", X"F9", X"9B", X"3E", X"BC", X"1F", X"FD", X"9E", 
        X"6E", X"6B", X"27", X"FD", X"9E", X"6E", X"6B", X"28", 
        X"00", X"A9", X"07", X"A0", X"E2", X"20", X"0E", X"E9", 
        X"A5", X"76", X"A6", X"75", X"85", X"9E", X"86", X"9F", 
        X"A2", X"90", X"38", X"20", X"45", X"F8", X"20", X"D4", 
        X"F9", X"4C", X"0E", X"E9", X"A0", X"01", X"A9", X"2D", 
        X"88", X"24", X"A2", X"10", X"04", X"C8", X"99", X"FF", 
        X"00", X"85", X"A2", X"84", X"AD", X"C8", X"A9", X"30", 
        X"A6", X"9D", X"D0", X"03", X"4C", X"F7", X"FA", X"A9", 
        X"00", X"E0", X"80", X"F0", X"02", X"B0", X"09", X"A9", 
        X"B4", X"A0", X"F9", X"20", X"29", X"F6", X"A9", X"F7", 
        X"85", X"99", X"A9", X"AF", X"A0", X"F9", X"20", X"57", 
        X"F8", X"F0", X"1E", X"10", X"12", X"A9", X"AA", X"A0", 
        X"F9", X"20", X"57", X"F8", X"F0", X"02", X"10", X"0E", 
        X"20", X"DE", X"F6", X"C6", X"99", X"D0", X"EE", X"20", 
        X"FA", X"F6", X"E6", X"99", X"D0", X"DC", X"20", X"4A", 
        X"F4", X"20", X"94", X"F8", X"A2", X"01", X"A5", X"99", 
        X"18", X"69", X"0A", X"30", X"09", X"C9", X"0B", X"B0", 
        X"06", X"69", X"FF", X"AA", X"A9", X"02", X"38", X"E9", 
        X"02", X"85", X"9A", X"86", X"99", X"8A", X"F0", X"02", 
        X"10", X"13", X"A4", X"AD", X"A9", X"2E", X"C8", X"99", 
        X"FF", X"00", X"8A", X"F0", X"06", X"A9", X"30", X"C8", 
        X"99", X"FF", X"00", X"84", X"AD", X"A0", X"00", X"A2", 
        X"80", X"A5", X"A1", X"18", X"79", X"0C", X"FB", X"85", 
        X"A1", X"A5", X"A0", X"79", X"0B", X"FB", X"85", X"A0", 
        X"A5", X"9F", X"79", X"0A", X"FB", X"85", X"9F", X"A5", 
        X"9E", X"79", X"09", X"FB", X"85", X"9E", X"E8", X"B0", 
        X"04", X"10", X"DE", X"30", X"02", X"30", X"DA", X"8A", 
        X"90", X"04", X"49", X"FF", X"69", X"0A", X"69", X"2F", 
        X"C8", X"C8", X"C8", X"C8", X"84", X"83", X"A4", X"AD", 
        X"C8", X"AA", X"29", X"7F", X"99", X"FF", X"00", X"C6", 
        X"99", X"D0", X"06", X"A9", X"2E", X"C8", X"99", X"FF", 
        X"00", X"84", X"AD", X"A4", X"83", X"8A", X"49", X"FF", 
        X"29", X"80", X"AA", X"C0", X"24", X"D0", X"AA", X"A4", 
        X"AD", X"B9", X"FF", X"00", X"88", X"C9", X"30", X"F0", 
        X"F8", X"C9", X"2E", X"F0", X"01", X"C8", X"A9", X"2B", 
        X"A6", X"9A", X"F0", X"2E", X"10", X"08", X"A9", X"00", 
        X"38", X"E5", X"9A", X"AA", X"A9", X"2D", X"99", X"01", 
        X"01", X"A9", X"45", X"99", X"00", X"01", X"8A", X"A2", 
        X"2F", X"38", X"E8", X"E9", X"0A", X"B0", X"FB", X"69", 
        X"3A", X"99", X"03", X"01", X"8A", X"99", X"02", X"01", 
        X"A9", X"00", X"99", X"04", X"01", X"F0", X"08", X"99", 
        X"FF", X"00", X"A9", X"00", X"99", X"00", X"01", X"A9", 
        X"00", X"A0", X"01", X"60", X"80", X"00", X"00", X"00", 
        X"00", X"FA", X"0A", X"1F", X"00", X"00", X"98", X"96", 
        X"80", X"FF", X"F0", X"BD", X"C0", X"00", X"01", X"86", 
        X"A0", X"FF", X"FF", X"D8", X"F0", X"00", X"00", X"03", 
        X"E8", X"FF", X"FF", X"FF", X"9C", X"00", X"00", X"00", 
        X"0A", X"FF", X"FF", X"FF", X"FF", X"20", X"08", X"F8", 
        X"A9", X"04", X"A0", X"FB", X"20", X"9E", X"F7", X"F0", 
        X"6F", X"A5", X"A5", X"D0", X"03", X"4C", X"FA", X"F4", 
        X"A2", X"8A", X"A0", X"00", X"20", X"D0", X"F7", X"A5", 
        X"AA", X"10", X"0F", X"20", X"C5", X"F8", X"A9", X"8A", 
        X"A0", X"00", X"20", X"57", X"F8", X"D0", X"03", X"98", 
        X"A4", X"0D", X"20", X"FA", X"F7", X"98", X"48", X"20", 
        X"EB", X"F5", X"A9", X"8A", X"A0", X"00", X"20", X"29", 
        X"F6", X"20", X"A8", X"FB", X"68", X"10", X"0A", X"A5", 
        X"9D", X"F0", X"06", X"A5", X"A2", X"49", X"FF", X"85", 
        X"A2", X"60", X"81", X"38", X"AA", X"3B", X"29", X"07", 
        X"71", X"34", X"58", X"3E", X"56", X"74", X"16", X"7E", 
        X"B3", X"1B", X"77", X"2F", X"EE", X"E3", X"85", X"7A", 
        X"1D", X"84", X"1C", X"2A", X"7C", X"63", X"59", X"58", 
        X"0A", X"7E", X"75", X"FD", X"E7", X"C6", X"80", X"31", 
        X"72", X"18", X"10", X"81", X"00", X"00", X"00", X"00", 
        X"A9", X"7A", X"A0", X"FB", X"20", X"29", X"F6", X"A5", 
        X"AC", X"69", X"50", X"90", X"03", X"20", X"1F", X"F8", 
        X"85", X"92", X"20", X"0B", X"F8", X"A5", X"9D", X"C9", 
        X"88", X"90", X"03", X"20", X"D0", X"F6", X"20", X"C5", 
        X"F8", X"A5", X"0D", X"18", X"69", X"81", X"F0", X"F3", 
        X"38", X"E9", X"01", X"48", X"A2", X"05", X"B5", X"A5", 
        X"B4", X"9D", X"95", X"9D", X"94", X"A5", X"CA", X"10", 
        X"F5", X"A5", X"92", X"85", X"AC", X"20", X"54", X"F4", 
        X"20", X"6F", X"FB", X"A9", X"7F", X"A0", X"FB", X"20", 
        X"10", X"FC", X"A9", X"00", X"85", X"AB", X"68", X"4C", 
        X"B8", X"F6", X"85", X"AD", X"84", X"AE", X"20", X"C6", 
        X"F7", X"A9", X"93", X"20", X"29", X"F6", X"20", X"14", 
        X"FC", X"A9", X"93", X"A0", X"00", X"4C", X"29", X"F6", 
        X"85", X"AD", X"84", X"AE", X"20", X"C3", X"F7", X"B1", 
        X"AD", X"85", X"A3", X"A4", X"AD", X"C8", X"98", X"D0", 
        X"02", X"E6", X"AE", X"85", X"AD", X"A4", X"AE", X"20", 
        X"29", X"F6", X"A5", X"AD", X"A4", X"AE", X"18", X"69", 
        X"05", X"90", X"01", X"C8", X"85", X"AD", X"84", X"AE", 
        X"20", X"68", X"F4", X"A9", X"98", X"A0", X"00", X"C6", 
        X"A3", X"D0", X"E4", X"60", X"98", X"35", X"44", X"7A", 
        X"68", X"28", X"B1", X"46", X"20", X"27", X"F8", X"AA", 
        X"30", X"18", X"A9", X"C9", X"A0", X"00", X"20", X"9E", 
        X"F7", X"8A", X"F0", X"E7", X"A9", X"44", X"A0", X"FC", 
        X"20", X"29", X"F6", X"A9", X"48", X"A0", X"FC", X"20", 
        X"68", X"F4", X"A6", X"A1", X"A5", X"9E", X"85", X"A1", 
        X"86", X"9E", X"A9", X"00", X"85", X"A2", X"A5", X"9D", 
        X"85", X"AC", X"A9", X"80", X"85", X"9D", X"20", X"D8", 
        X"F4", X"A2", X"C9", X"A0", X"00", X"4C", X"D0", X"F7", 
        X"E6", X"B8", X"D0", X"02", X"E6", X"B9", X"AD", X"60", 
        X"EA", X"C9", X"3A", X"B0", X"0A", X"C9", X"20", X"F0", 
        X"EF", X"38", X"E9", X"30", X"38", X"E9", X"D0", X"60", 
        X"80", X"4F", X"C7", X"52", X"58", X"A2", X"FF", X"86", 
        X"76", X"A2", X"FB", X"9A", X"A9", X"A5", X"A0", X"FC", 
        X"85", X"01", X"84", X"02", X"85", X"04", X"84", X"05", 
        X"A9", X"4C", X"85", X"00", X"85", X"03", X"85", X"90", 
        X"A2", X"1C", X"BD", X"87", X"FC", X"95", X"B0", X"CA", 
        X"D0", X"F8", X"8A", X"85", X"A4", X"85", X"54", X"48", 
        X"A9", X"03", X"85", X"8F", X"20", X"34", X"FE", X"A9", 
        X"01", X"8D", X"FD", X"01", X"8D", X"FC", X"01", X"A2", 
        X"55", X"86", X"52", X"A9", X"00", X"A0", X"08", X"85", 
        X"50", X"84", X"51", X"A0", X"00", X"E6", X"51", X"B1", 
        X"50", X"49", X"FF", X"91", X"50", X"D1", X"50", X"D0", 
        X"08", X"49", X"FF", X"91", X"50", X"D1", X"50", X"F0", 
        X"EC", X"A4", X"50", X"A5", X"51", X"29", X"F0", X"84", 
        X"73", X"85", X"74", X"84", X"6F", X"85", X"70", X"A2", 
        X"00", X"A0", X"08", X"86", X"67", X"84", X"68", X"A0", 
        X"00", X"84", X"D6", X"98", X"91", X"67", X"E6", X"67", 
        X"D0", X"02", X"E6", X"68", X"A5", X"67", X"A4", X"68", 
        X"20", X"91", X"E2", X"20", X"D2", X"E4", X"A9", X"0E", 
        X"A0", X"E9", X"85", X"04", X"84", X"05", X"A9", X"EA", 
        X"A0", X"E2", X"85", X"01", X"84", X"02", X"6C", X"01", 
        X"00", X"20", X"17", X"EB", X"20", X"18", X"F4", X"6C", 
        X"50", X"00", X"20", X"17", X"EB", X"20", X"18", X"F4", 
        X"A5", X"50", X"C5", X"6D", X"A5", X"51", X"E5", X"6E", 
        X"B0", X"03", X"4C", X"BE", X"E2", X"A5", X"50", X"85", 
        X"73", X"85", X"6F", X"A5", X"51", X"85", X"74", X"85", 
        X"70", X"60", X"20", X"17", X"EB", X"20", X"18", X"F4", 
        X"A5", X"50", X"C5", X"73", X"A5", X"51", X"E5", X"74", 
        X"B0", X"E0", X"A5", X"50", X"C5", X"69", X"A5", X"51", 
        X"E5", X"6A", X"90", X"D6", X"A5", X"50", X"85", X"69", 
        X"A5", X"51", X"85", X"6A", X"4C", X"F3", X"E4", X"A9", 
        X"8E", X"20", X"69", X"EC", X"A5", X"B8", X"85", X"F4", 
        X"A5", X"B9", X"85", X"F5", X"38", X"66", X"D8", X"A5", 
        X"75", X"85", X"F6", X"A5", X"76", X"85", X"F7", X"20", 
        X"A2", X"E7", X"4C", X"94", X"E7", X"86", X"DE", X"A6", 
        X"F8", X"86", X"DF", X"A5", X"75", X"85", X"DA", X"A5", 
        X"76", X"85", X"DB", X"A5", X"79", X"85", X"DC", X"A5", 
        X"7A", X"85", X"DD", X"A5", X"F4", X"85", X"B8", X"A5", 
        X"F5", X"85", X"B9", X"A5", X"F6", X"85", X"75", X"A5", 
        X"F7", X"85", X"76", X"20", X"B7", X"00", X"20", X"3A", 
        X"E7", X"4C", X"48", X"E6", X"A5", X"DA", X"85", X"75", 
        X"A5", X"DB", X"85", X"76", X"A5", X"DC", X"85", X"B8", 
        X"A5", X"DD", X"85", X"B9", X"A6", X"DF", X"9A", X"4C", 
        X"48", X"E6", X"AD", X"11", X"D0", X"10", X"FB", X"AD", 
        X"10", X"D0", X"29", X"7F", X"60", X"C9", X"18", X"F0", 
        X"0A", X"20", X"EF", X"FF", X"C9", X"5F", X"F0", X"0E", 
        X"E8", X"D0", X"0F", X"20", X"28", X"FE", X"20", X"34", 
        X"FE", X"20", X"2B", X"FE", X"A2", X"01", X"8A", X"F0", 
        X"F5", X"CA", X"20", X"F2", X"FD", X"9D", X"00", X"02", 
        X"C9", X"0D", X"D0", X"D9", X"20", X"34", X"FE", X"60", 
        X"A9", X"5C", X"2C", X"A5", X"33", X"2C", X"A9", X"20", 
        X"2C", X"A9", X"3F", X"2C", X"A9", X"0D", X"09", X"80", 
        X"20", X"EF", X"FF", X"29", X"7F", X"60", X"A0", X"18", 
        X"20", X"34", X"FE", X"88", X"10", X"FA", X"60", X"AC", 
        X"DC", X"AF", X"C0", X"CF", X"D0", X"5B", X"AC", X"DD", 
        X"AF", X"C0", X"FA", X"D0", X"54", X"60", X"20", X"47", 
        X"FE", X"4C", X"06", X"90", X"20", X"47", X"FE", X"A0", 
        X"00", X"B9", X"00", X"00", X"99", X"80", X"03", X"C8", 
        X"C0", X"0C", X"D0", X"F5", X"C6", X"B8", X"A0", X"00", 
        X"20", X"B1", X"00", X"F0", X"08", X"99", X"C1", X"03", 
        X"C8", X"C0", X"0F", X"D0", X"F3", X"C0", X"00", X"F0", 
        X"2B", X"8C", X"C0", X"03", X"A9", X"C0", X"A0", X"03", 
        X"85", X"02", X"84", X"03", X"A5", X"AF", X"E5", X"67", 
        X"85", X"09", X"A5", X"B0", X"E5", X"68", X"85", X"0A", 
        X"A5", X"67", X"A4", X"68", X"85", X"00", X"85", X"07", 
        X"84", X"01", X"84", X"08", X"A9", X"F8", X"85", X"06", 
        X"60", X"A2", X"8C", X"2C", X"A2", X"06", X"4C", X"C0", 
        X"E2", X"A0", X"00", X"B9", X"80", X"03", X"99", X"00", 
        X"00", X"C8", X"C0", X"0C", X"D0", X"F5", X"60", X"20", 
        X"5C", X"FE", X"A2", X"20", X"20", X"E5", X"FE", X"20", 
        X"B1", X"FE", X"60", X"20", X"5C", X"FE", X"A2", X"22", 
        X"20", X"E5", X"FE", X"A5", X"67", X"65", X"09", X"85", 
        X"69", X"A5", X"68", X"65", X"0A", X"85", X"6A", X"20", 
        X"B1", X"FE", X"4C", X"A0", X"E3", X"20", X"0C", X"90", 
        X"A2", X"04", X"B0", X"F9", X"60", X"00", X"00", X"00", 
        X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
        X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
        X"D8", X"58", X"A0", X"7F", X"8C", X"12", X"D0", X"A9", 
        X"A7", X"8D", X"11", X"D0", X"8D", X"13", X"D0", X"C9", 
        X"DF", X"F0", X"13", X"C9", X"9B", X"F0", X"03", X"C8", 
        X"10", X"0F", X"A9", X"DC", X"20", X"EF", X"FF", X"A9", 
        X"8D", X"20", X"EF", X"FF", X"A0", X"01", X"88", X"30", 
        X"F6", X"AD", X"11", X"D0", X"10", X"FB", X"AD", X"10", 
        X"D0", X"99", X"00", X"02", X"20", X"EF", X"FF", X"C9", 
        X"8D", X"D0", X"D4", X"A0", X"FF", X"A9", X"00", X"AA", 
        X"0A", X"85", X"2B", X"C8", X"B9", X"00", X"02", X"C9", 
        X"8D", X"F0", X"D4", X"C9", X"AE", X"90", X"F4", X"F0", 
        X"F0", X"C9", X"BA", X"F0", X"EB", X"C9", X"D2", X"F0", 
        X"3B", X"86", X"28", X"86", X"29", X"84", X"2A", X"B9", 
        X"00", X"02", X"49", X"B0", X"C9", X"0A", X"90", X"06", 
        X"69", X"88", X"C9", X"FA", X"90", X"11", X"0A", X"0A", 
        X"0A", X"0A", X"A2", X"04", X"0A", X"26", X"28", X"26", 
        X"29", X"CA", X"D0", X"F8", X"C8", X"D0", X"E0", X"C4", 
        X"2A", X"F0", X"97", X"24", X"2B", X"50", X"10", X"A5", 
        X"28", X"81", X"26", X"E6", X"26", X"D0", X"B5", X"E6", 
        X"27", X"4C", X"44", X"FF", X"6C", X"24", X"00", X"30", 
        X"2B", X"A2", X"02", X"B5", X"27", X"95", X"25", X"95", 
        X"23", X"CA", X"D0", X"F7", X"D0", X"14", X"A9", X"8D", 
        X"20", X"EF", X"FF", X"A5", X"25", X"20", X"DC", X"FF", 
        X"A5", X"24", X"20", X"DC", X"FF", X"A9", X"BA", X"20", 
        X"EF", X"FF", X"A9", X"A0", X"20", X"EF", X"FF", X"A1", 
        X"24", X"20", X"DC", X"FF", X"86", X"2B", X"A5", X"24", 
        X"C5", X"28", X"A5", X"25", X"E5", X"29", X"B0", X"C1", 
        X"E6", X"24", X"D0", X"02", X"E6", X"25", X"A5", X"24", 
        X"29", X"07", X"10", X"C8", X"48", X"4A", X"4A", X"4A", 
        X"4A", X"20", X"E5", X"FF", X"68", X"29", X"0F", X"09", 
        X"B0", X"C9", X"BA", X"90", X"02", X"69", X"06", X"2C", 
        X"12", X"D0", X"30", X"FB", X"8D", X"12", X"D0", X"60", 
        X"00", X"00", X"00", X"0F", X"00", X"FF", X"00", X"00"
    );
begin
    process(clock)
    begin
        if rising_edge(clock) then
            if cs_n = '0' then
                data_out <= rom(to_integer(unsigned(address)));
            end if;
        end if;
    end process;

end rtl;
