library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cpu_timing is
    generic (
        SDRAM_MHZ : integer := 100;  -- SDRAM clock frequency
        CPU_MHZ   : integer := 10    -- CPU (PHI2) frequency
    );
    port (
        clk       : in  std_logic;   -- SDRAM clock
        phi2      : in  std_logic;   -- CPU PHI2 input
        reset     : in  std_logic;
        
        -- Timing outputs
        phi2_early : out std_logic;  -- Early in PHI2 cycle
        phi2_mid   : out std_logic;  -- Middle of PHI2 cycle
        phi2_late  : out std_logic;  -- Late in PHI2 cycle (before fall)
        phi2_rise  : out std_logic;  -- Single-cycle pulse on PHI2 rising
        phi2_fall  : out std_logic   -- Single-cycle pulse on PHI2 falling
    );
end cpu_timing;

architecture rtl of cpu_timing is
    -- Calculate SDRAM cycles during PHI2 HIGH (assuming 50% duty cycle)
    constant PHI2_HIGH_NS : integer := (1000 / (2 * CPU_MHZ));
    constant SDRAM_CYCLES : integer := (SDRAM_MHZ * PHI2_HIGH_NS) / 1000;
    
    -- Define timing windows (in SDRAM cycles)
    constant EARLY_END : integer := 1;
    constant MID_END   : integer := SDRAM_CYCLES / 2;
    constant LATE_START : integer := SDRAM_CYCLES - 2;
    
    signal phi2_prev  : std_logic;
    signal phase_counter : integer range 0 to 63;
    
begin
    process(clk)
    begin
        if rising_edge(clk) then
            phi2_prev <= phi2;
            
            if reset = '1' then
                phase_counter <= 0;
                phi2_early <= '0';
                phi2_mid <= '0';
                phi2_late <= '0';
                phi2_rise <= '0';
                phi2_fall <= '0';
            else
                -- Detect edges
                phi2_rise <= '1' when (phi2 = '1' and phi2_prev = '0') else '0';
                phi2_fall <= '1' when (phi2 = '0' and phi2_prev = '1') else '0';
                
                -- Phase counter
                if phi2 = '1' and phi2_prev = '0' then
                    phase_counter <= 0;
                elsif phi2 = '1' then
                    if phase_counter < 63 then
                        phase_counter <= phase_counter + 1;
                    end if;
                end if;
                
                -- Generate timing windows
                phi2_early <= '1' when (phi2 = '1' and phase_counter <= EARLY_END) else '0';
                phi2_mid   <= '1' when (phi2 = '1' and phase_counter > EARLY_END and phase_counter < LATE_START) else '0';
                phi2_late  <= '1' when (phi2 = '1' and phase_counter >= LATE_START) else '0';
            end if;
        end if;
    end process;
    
end rtl;