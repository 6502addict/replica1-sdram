-- Simple SDRAM Controller Template for Logic Analyzer Debug
-- 100MHz operation for IS42S16320F
-- Write your own logic from here!

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sdram_controller is
    generic (
	     FREQ_MHZ : integer := 100; -- Clock frequency in MHz
        ROW_BITS : integer := 13;  -- 13 for DE10-Lite, 12 for DE1
        COL_BITS : integer := 10   -- 10 for DE10-Lite, 8 for DE1
    );
    port(
        clk         : in    std_logic;  -- 20MHz
        reset       : in    std_logic;  -- Active high
        
        -- Simple CPU interface
        req         : in    std_logic;
        wr          : in    std_logic;  -- 1=write, 0=read
		  addr        : in    std_logic_vector(ROW_BITS+COL_BITS+1 downto 0); 
        din         : in    std_logic_vector(15 downto 0);
        dout        : out   std_logic_vector(15 downto 0);
        byte_en     : in    std_logic_vector(1 downto 0);  -- Active low (not used yet, always "00")
        ready       : out   std_logic;
        ack         : out   std_logic;
        
        -- Debug outputs for logic analyzer
        debug_state    : out   std_logic_vector(3 downto 0);  -- Current FSM state
        debug_cmd      : out   std_logic_vector(3 downto 0);  -- Current SDRAM command
--      debug_seq      : out   std_logic_vector(15 downto 0);  -- Sequence counter (lower 8 bits)
        refresh_active : out   std_logic;  -- High during refresh
        
        -- SDRAM pins
        sdram_clk   : out   std_logic;
        sdram_cke   : out   std_logic;
        sdram_cs_n  : out   std_logic;
        sdram_ras_n : out   std_logic;
        sdram_cas_n : out   std_logic;
        sdram_we_n  : out   std_logic;
        sdram_ba    : out   std_logic_vector(1 downto 0);
        sdram_addr  : out   std_logic_vector(12 downto 0);
        sdram_dq    : inout std_logic_vector(15 downto 0);
        sdram_dqm   : out   std_logic_vector(1 downto 0)
    );
end sdram_controller;

architecture rtl of sdram_controller is

    -- SDRAM Commands (CS_N, RAS_N, CAS_N, WE_N)
    constant CMD_NOP       : std_logic_vector(3 downto 0) := "0111";
    constant CMD_ACTIVE    : std_logic_vector(3 downto 0) := "0011";
    constant CMD_READ      : std_logic_vector(3 downto 0) := "0101";
    constant CMD_WRITE     : std_logic_vector(3 downto 0) := "0100";
    constant CMD_PRECHARGE : std_logic_vector(3 downto 0) := "0010";
    constant CMD_REFRESH   : std_logic_vector(3 downto 0) := "0001";
    constant CMD_LOAD_MODE : std_logic_vector(3 downto 0) := "0000";
    
    -- States (visible on logic analyzer via debug_state)
    constant ST_INIT       : std_logic_vector(3 downto 0) := "0000";
    constant ST_IDLE       : std_logic_vector(3 downto 0) := "0001";
    constant ST_REFRESH    : std_logic_vector(3 downto 0) := "0010";
    constant ST_ACTIVATE   : std_logic_vector(3 downto 0) := "0011";
    constant ST_READ       : std_logic_vector(3 downto 0) := "0100";
    constant ST_WRITE      : std_logic_vector(3 downto 0) := "0101";
    constant ST_PRECHARGE  : std_logic_vector(3 downto 0) := "0110";
	 
	 -- SDRAM timing parameters (in nanoseconds)
  	 constant TRP_NS  : integer := 20;   -- Precharge time
	 constant TRCD_NS : integer := 20;   -- RAS to CAS delay
	 constant TRFC_NS : integer := 70;   -- Refresh cycle time

	 -- Compute cycles needed (round up)
	 constant TRP_CYCLES  : integer := ((TRP_NS * FREQ_MHZ) + 999) / 1000;
	 constant TRCD_CYCLES : integer := ((TRCD_NS * FREQ_MHZ) + 999) / 1000;
	 constant TRFC_CYCLES : integer := ((TRFC_NS * FREQ_MHZ) + 999) / 1000;

 	 constant INIT_WAIT        : integer := FREQ_MHZ * 200;      -- 200µs
	 constant REFRESH_INTERVAL : integer := (FREQ_MHZ * 78) / 10; -- 7.8µs

    signal state : std_logic_vector(3 downto 0) := ST_INIT;
	 signal seq_count : integer range 0 to INIT_WAIT + 50 := 0;

    
    signal refresh_counter : integer range 0 to REFRESH_INTERVAL := 0;
    signal need_refresh : std_logic := '0';
    signal init_done : std_logic := '0';  -- Flag: initialization complete
    
    -- Command outputs
    signal cmd : std_logic_vector(3 downto 0) := CMD_NOP;
    
    -- Address latches
    signal addr_bank : std_logic_vector(1 downto 0);
    signal addr_row  : std_logic_vector(ROW_BITS-1 downto 0);
    signal addr_col  : std_logic_vector(COL_BITS-1 downto 0);
    signal data_out  : std_logic_vector(15 downto 0);
	 
	 signal sdram_cs_n_reg  : std_logic;
    signal sdram_ras_n_reg : std_logic;
    signal sdram_cas_n_reg : std_logic;
    signal sdram_we_n_reg  : std_logic;
    signal sdram_ba_reg    : std_logic_vector(1 downto 0);
    signal sdram_addr_reg  : std_logic_vector(12 downto 0);
    signal sdram_dqm_reg   : std_logic_vector(1 downto 0);

begin

    -- Output assignments
    sdram_clk <= clk;
    sdram_cke <= '1';
    sdram_cs_n  <= sdram_cs_n_reg;
    sdram_ras_n <= sdram_ras_n_reg;
    sdram_cas_n <= sdram_cas_n_reg;
    sdram_we_n  <= sdram_we_n_reg;
    sdram_ba    <= sdram_ba_reg;
    sdram_addr  <= sdram_addr_reg;
    sdram_dqm   <= sdram_dqm_reg;	 
--    sdram_cs_n  <= cmd(3);
--    sdram_ras_n <= cmd(2);
--    sdram_cas_n <= cmd(1);
--    sdram_we_n  <= cmd(0);
    
    -- Debug outputs
    debug_state <= state;
    debug_cmd <= cmd;  -- Show command being sent
--    debug_seq <= std_logic_vector(to_unsigned(seq_count, 16));  -- 16 bits of counter
    refresh_active <= '1' when state = ST_REFRESH else '0';
    
    -- Data bus (tristate when not writing)
    sdram_dq <= din when (state = ST_WRITE and seq_count = 0) else (others => 'Z');
    
    process(clk)
    begin
        if rising_edge(clk) then
            sdram_cs_n_reg  <= cmd(3);
            sdram_ras_n_reg <= cmd(2);
            sdram_cas_n_reg <= cmd(1);
            sdram_we_n_reg  <= cmd(0);		  
		  
            if reset = '1' then
                state <= ST_INIT;
                seq_count <= 0;
                cmd <= CMD_NOP;
                sdram_ba_reg <= "00";
                sdram_addr_reg <= (others => '0');
                sdram_dqm_reg <= "11";
                ready <= '0';
                ack <= '0';
                refresh_counter <= 0;
                need_refresh <= '0';
                init_done <= '0';
                
            else
                -- Default: clear ack
                ack <= '0';
                
                -- Refresh counter (ONLY after initialization complete)
                if init_done = '1' then
                    if refresh_counter >= REFRESH_INTERVAL then
                        refresh_counter <= 0;
                        need_refresh <= '1';
                    else
                        refresh_counter <= refresh_counter + 1;
                    end if;
                end if;
                
                case state is
                    
                    --========================================
                    -- INITIALIZATION
                    --========================================
                    when ST_INIT =>
                        ready <= '0';
                        cmd <= CMD_NOP;
                        
                        if seq_count < INIT_WAIT then
                            -- Wait 200us
                            seq_count <= seq_count + 1;
                            
                        elsif seq_count = INIT_WAIT then
                            -- PRECHARGE ALL
                            cmd <= CMD_PRECHARGE;
                            sdram_addr_reg(10) <= '1';  -- All banks
                            seq_count <= seq_count + 1;
                            
                        elsif seq_count = INIT_WAIT + 2 then
                            -- First REFRESH
                            cmd <= CMD_REFRESH;
                            seq_count <= seq_count + 1;
                            
                        elsif seq_count = INIT_WAIT + 10 then
                            -- Second REFRESH
                            cmd <= CMD_REFRESH;
                            seq_count <= seq_count + 1;
                            
                        elsif seq_count = INIT_WAIT + 18 then
                            -- MODE REGISTER SET
                            -- CAS=2, Sequential, Burst=1
                            cmd <= CMD_LOAD_MODE;
                            sdram_ba_reg <= "00";
                            sdram_addr_reg <= "0000" & "00" & "010" & "0" & "000";
                            seq_count <= seq_count + 1;
                            
                        elsif seq_count = INIT_WAIT + 20 then
                            -- Done! Go to IDLE
                            cmd <= CMD_NOP;
                            state <= ST_IDLE;
                            seq_count <= 0;
                            ready <= '1';
                            init_done <= '1';  -- Enable refresh counter
                            
                        else
                            cmd <= CMD_NOP;
                            seq_count <= seq_count + 1;
                        end if;
                    
                    --========================================
                    -- IDLE - Wait for request or refresh
                    --========================================
                    when ST_IDLE =>
                        cmd <= CMD_NOP;
                        sdram_dqm_reg <= "11";
                        ready <= '1';
                        seq_count <= 0;
                        
                        if need_refresh = '1' then
                            -- Do refresh
                            state <= ST_REFRESH;
                            ready <= '0';
                            
                        elsif req = '1' then
                            -- Latch address
                            addr_bank <= addr(addr'high downto addr'high-1);
                            addr_row <= addr(addr'high-2 downto COL_BITS);
                            addr_col <= addr(COL_BITS-1 downto 0);
                            state <= ST_ACTIVATE;
                            ready <= '0';
                        end if;
                    
                    --========================================
                    -- REFRESH
                    --========================================
                    when ST_REFRESH =>
                        if seq_count = 0 then
                            cmd <= CMD_REFRESH;
                            seq_count <= seq_count + 1;
                        elsif seq_count = TRFC_CYCLES then
                            cmd <= CMD_NOP;
                            need_refresh <= '0';
                            state <= ST_IDLE;
                            seq_count <= 0;
                        else
                            cmd <= CMD_NOP;
                            seq_count <= seq_count + 1;
                        end if;
                    
                    --========================================
                    -- ACTIVATE ROW
                    --========================================
                    when ST_ACTIVATE =>
                        if seq_count = 0 then
                            cmd <= CMD_ACTIVE;
                            sdram_ba_reg <= addr_bank;
									 sdram_addr_reg <= std_logic_vector(resize(unsigned(addr_row), 13));
                            seq_count <= seq_count + 1;
                        elsif seq_count = TRCD_CYCLES then
                            cmd <= CMD_NOP;
                            -- Decide read or write
                            if wr = '1' then
                                state <= ST_WRITE;
                            else
                                state <= ST_READ;
                            end if;
                            seq_count <= 0;
                        else
                            cmd <= CMD_NOP;
                            seq_count <= seq_count + 1;
                        end if;
                    
                    --========================================
                    -- READ
                    --========================================
                    when ST_READ =>
                        if seq_count = 0 then
                            -- Issue READ command with auto-precharge
                            cmd <= CMD_READ;
                            sdram_ba_reg <= addr_bank;
									 sdram_addr_reg <= (others => '0');
									 sdram_addr_reg(10) <= '1';  -- A10=1 for auto-precharge
									 sdram_addr_reg(COL_BITS-1 downto 0) <= addr_col;
									 sdram_dqm_reg <= not byte_en;
                            seq_count <= seq_count + 1;
                            
                        elsif seq_count = TRP_CYCLES then
                            -- Data available (CAS latency = 2)
                            cmd <= CMD_NOP;
                            dout <= sdram_dq;
                            ack <= '1';
                            sdram_dqm_reg <= "11";
                            seq_count <= seq_count + 1;
                            
                        elsif seq_count = 5 then
                            -- Auto-precharge complete, back to idle
                            state <= ST_IDLE;
                            seq_count <= 0;
                            
                        else
                            cmd <= CMD_NOP;
                            seq_count <= seq_count + 1;
                        end if;
                    
                    --========================================
                    -- WRITE
                    --========================================
                    when ST_WRITE =>
                        if seq_count = 0 then
                            -- Issue WRITE command with auto-precharge
                            cmd <= CMD_WRITE;
                            sdram_ba_reg <= addr_bank;
									 sdram_addr_reg <= (others => '0');
									 sdram_addr_reg(10) <= '1';  -- A10=1 for auto-precharge
								    sdram_addr_reg(COL_BITS-1 downto 0) <= addr_col;
									 sdram_dqm_reg <= not byte_en;
                            -- din is on data bus (see concurrent assignment)
                            ack <= '1';
                            seq_count <= seq_count + 1;
                            
                        elsif seq_count = TRP_CYCLES then
                            -- Auto-precharge complete, back to idle
                            cmd <= CMD_NOP;
                            sdram_dqm_reg <= "11";
                            state <= ST_IDLE;
                            seq_count <= 0;
                            
                        else
                            cmd <= CMD_NOP;
                            seq_count <= seq_count + 1;
                        end if;
                    
                    when others =>
                        state <= ST_INIT;
                        
                end case;
            end if;
        end if;
    end process;

end rtl;