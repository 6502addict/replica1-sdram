-- ============================================================================
-- Apple1_CPU_6800.vhd
-- Derived from Apple1_CPU_Template.vhd
-- 
-- CPU: MC6800 (Motorola 6800 8-bit processor)
-- Dependencies: None (uses standard IEEE libraries only)
-- Note: This creates a "6800-based Apple 1" - different instruction set!
-- https://opencores.org/projects/system68
-- ============================================================================

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity CPU_6800 is
	port (
		-- Clock and Reset
		main_clk : in  std_logic;       -- Main system clock
		reset_n  : in  std_logic;       -- Active low reset
		phi2     : out std_logic;       -- Phase 2 clock output (divided from main_clk)
		
		-- CPU Control Interface
		rw       : out std_logic;       -- Read/Write (1=Read, 0=Write)
		vma      : out std_logic;       -- Valid Memory Access
		sync     : out std_logic;       -- Instruction fetch cycle
		
		-- Address and Data Bus
		addr     : out std_logic_vector(15 downto 0);  -- Address bus
		data_in  : in  std_logic_vector(7 downto 0);   -- Data input
		data_out : out std_logic_vector(7 downto 0);   -- Data output
		
		-- Interrupt Interface  
		nmi_n    : in  std_logic;       -- Non-maskable interrupt (active low)
		irq_n    : in  std_logic;       -- Interrupt request (active low)
		so_n     : in  std_logic := '1' -- Set overflow (not used by 6800)
	);
end CPU_6800;

architecture MC6800_impl of CPU_6800 is


	component clock_divider is
		 generic (divider : integer := 4);
		 port (
			  reset    : in  std_logic := '1';
			  clk_in   : in  std_logic;
			  clk_out  : out std_logic
		 );
	end component;

	-- MC6800 Component (cpu68 core)
	component cpu68 is
		port (
			clk     : in std_logic;                         -- Clock (main_clk)
			rst     : in std_logic;                         -- Reset (active high)
			rw      : out std_logic;                        -- Read/Write
			vma     : out std_logic;                        -- Valid Memory Access
			address : out std_logic_vector(15 downto 0);    -- Address bus
			data_in : in std_logic_vector(7 downto 0);      -- Data input
			data_out: out std_logic_vector(7 downto 0);     -- Data output
			irq     : in std_logic;                         -- IRQ (active high)
			nmi     : in std_logic;                         -- NMI (active high)
			halt    : in std_logic;                         -- Halt
			hold    : in std_logic                          -- Hold/DMA request
		);
	end component;

	-- Internal signals
	signal reset_internal: std_logic;              -- Internal reset (active high)
	signal data_bus      : std_logic_vector(7 downto 0);
	signal address_bus   : std_logic_vector(15 downto 0);
	signal cpu_data_out  : std_logic_vector(7 downto 0);
	signal rw_internal   : std_logic;
	signal sync_internal : std_logic;
	signal vma_internal  : std_logic;
	signal phi2_internal : std_logic;

	-- MC6800 specific signals
	signal mc6800_rw     : std_logic;
	signal mc6800_vma    : std_logic;

begin

	clk:  clock_divider generic map(divider         => 2)  
								  port map(reset           => '1',
									  	     clk_in          => main_clk,
											  clk_out         => phi2_internal);	
											  
	phi2 <= phi2_internal;

	-- Clock and reset assignments
	reset_internal <= not reset_n;

	-- Input data bus assignment
	data_bus <= data_in;

	-- MC6800 Instantiation
	mc6800_inst: cpu68 
		port map(
			clk     => phi2_internal,              -- CPU68 uses main_clk directly
			rst     => reset_internal,             -- MC6800 uses active high reset
			rw      => mc6800_rw,
			vma     => mc6800_vma,
			address => address_bus,
			data_in => data_bus,
			data_out=> cpu_data_out,
			irq     => not irq_n,                  -- MC6800 uses active high
			nmi     => not nmi_n,                  -- MC6800 uses active high
			halt    => '0',                        -- No halt for Apple 1
			hold    => '0'                         -- No DMA for Apple 1
		);
		
	-- Signal assignments for MC6800
	rw_internal   <= mc6800_rw;
	vma_internal  <= mc6800_vma;                  -- MC6800 provides its own VMA
	sync_internal <= '0';                         -- 6800 doesn't have sync like 6502
	
	-- Note: 6800 VMA timing is different from 6502:
	-- - 6502: VMA = phi2 (address valid during phi2 high)
	-- - 6800: VMA is generated by CPU based on internal state

	-- Output assignments
	addr     <= address_bus;
	data_out <= cpu_data_out;
	rw       <= rw_internal;
	sync     <= sync_internal;
	vma      <= vma_internal;

end MC6800_impl;